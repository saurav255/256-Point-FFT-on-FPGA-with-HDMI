`timescale 1ns / 1ps

// This version is 8 point fft using ram 


module fft_ver2 #(
    parameter WIDTH = 20  // bit-width for fixed-point
)(input clk, rst, trig, input [((2*WIDTH)-1):0]doutb, input [((2*WIDTH)-1):0]dout_tw, output reg [((2*WIDTH)-1):0]douta, output reg [10:0]addr_tw, 
  output reg [7:0]addrb, output reg [7:0]addra, output reg wr, output reg done, output reg [23:0]d_fifo_ram, output reg wr_fifo_ram, 
  output reg [9:0]addr_fifo_ram, output [3:0]state_fft

    ); 
    
    localparam SHIFT_FACTOR = 8;
    
    // twiddle factor rom signals 
    reg [((2*WIDTH)-1):0]tw;

    
    // signal declarations for unit fft component  
    reg signed [WIDTH-1:0]in1_real;
    reg signed [WIDTH-1:0]in1_imag;
    reg signed [WIDTH-1:0]in2_real;
    reg signed [WIDTH-1:0]in2_imag;
    reg signed [WIDTH-1:0]w_real;
    reg signed [WIDTH-1:0]w_imag;
    wire signed [WIDTH-1:0]out1_real;
    wire signed [WIDTH-1:0]out1_imag;
    wire signed [WIDTH-1:0]out2_real;
    wire signed [WIDTH-1:0]out2_imag;
    
    // Unit instance 
    unit unit_1(
    // complex inputs
    .in1_real(in1_real),
    .in1_imag(in1_imag),
    .in2_real(in2_real),
    .in2_imag(in2_imag),

    // complex twiddle factor
    .w_real(w_real),
    .w_imag(w_imag),

    // complex outputs
    .out1_real(out1_real),
    .out1_imag(out1_imag),
    .out2_real(out2_real),
    .out2_imag(out2_imag)
    );
    // ====================== Index store =================
    reg [7:0]STAGE1_IND[0:255]; 
    reg [7:0]STAGE2_IND[0:255]; 
    reg [7:0]STAGE3_IND[0:255]; 
    reg [7:0]STAGE4_IND[0:255]; 
    reg [7:0]STAGE5_IND[0:255]; 
    reg [7:0]STAGE6_IND[0:255]; 
    reg [7:0]STAGE7_IND[0:255]; 
    reg [7:0]STAGE8_IND[0:255];
    reg [7:0]BITFLIP_IND[0:255]; 
initial begin
   STAGE1_IND[0] <= 8'd0;
    STAGE1_IND[1] <= 8'd128;
    STAGE1_IND[2] <= 8'd64;
    STAGE1_IND[3] <= 8'd192;
    STAGE1_IND[4] <= 8'd32;
    STAGE1_IND[5] <= 8'd160;
    STAGE1_IND[6] <= 8'd96;
    STAGE1_IND[7] <= 8'd224;
    STAGE1_IND[8] <= 8'd16;
    STAGE1_IND[9] <= 8'd144;
    STAGE1_IND[10] <= 8'd80;
    STAGE1_IND[11] <= 8'd208;
    STAGE1_IND[12] <= 8'd48;
    STAGE1_IND[13] <= 8'd176;
    STAGE1_IND[14] <= 8'd112;
    STAGE1_IND[15] <= 8'd240;
    STAGE1_IND[16] <= 8'd8;
    STAGE1_IND[17] <= 8'd136;
    STAGE1_IND[18] <= 8'd72;
    STAGE1_IND[19] <= 8'd200;
    STAGE1_IND[20] <= 8'd40;
    STAGE1_IND[21] <= 8'd168;
    STAGE1_IND[22] <= 8'd104;
    STAGE1_IND[23] <= 8'd232;
    STAGE1_IND[24] <= 8'd24;
    STAGE1_IND[25] <= 8'd152;
    STAGE1_IND[26] <= 8'd88;
    STAGE1_IND[27] <= 8'd216;
    STAGE1_IND[28] <= 8'd56;
    STAGE1_IND[29] <= 8'd184;
    STAGE1_IND[30] <= 8'd120;
    STAGE1_IND[31] <= 8'd248;
    STAGE1_IND[32] <= 8'd4;
    STAGE1_IND[33] <= 8'd132;
    STAGE1_IND[34] <= 8'd68;
    STAGE1_IND[35] <= 8'd196;
    STAGE1_IND[36] <= 8'd36;
    STAGE1_IND[37] <= 8'd164;
    STAGE1_IND[38] <= 8'd100;
    STAGE1_IND[39] <= 8'd228;
    STAGE1_IND[40] <= 8'd20;
    STAGE1_IND[41] <= 8'd148;
    STAGE1_IND[42] <= 8'd84;
    STAGE1_IND[43] <= 8'd212;
    STAGE1_IND[44] <= 8'd52;
    STAGE1_IND[45] <= 8'd180;
    STAGE1_IND[46] <= 8'd116;
    STAGE1_IND[47] <= 8'd244;
    STAGE1_IND[48] <= 8'd12;
    STAGE1_IND[49] <= 8'd140;
    STAGE1_IND[50] <= 8'd76;
    STAGE1_IND[51] <= 8'd204;
    STAGE1_IND[52] <= 8'd44;
    STAGE1_IND[53] <= 8'd172;
    STAGE1_IND[54] <= 8'd108;
    STAGE1_IND[55] <= 8'd236;
    STAGE1_IND[56] <= 8'd28;
    STAGE1_IND[57] <= 8'd156;
    STAGE1_IND[58] <= 8'd92;
    STAGE1_IND[59] <= 8'd220;
    STAGE1_IND[60] <= 8'd60;
    STAGE1_IND[61] <= 8'd188;
    STAGE1_IND[62] <= 8'd124;
    STAGE1_IND[63] <= 8'd252;
    STAGE1_IND[64] <= 8'd2;
    STAGE1_IND[65] <= 8'd130;
    STAGE1_IND[66] <= 8'd66;
    STAGE1_IND[67] <= 8'd194;
    STAGE1_IND[68] <= 8'd34;
    STAGE1_IND[69] <= 8'd162;
    STAGE1_IND[70] <= 8'd98;
    STAGE1_IND[71] <= 8'd226;
    STAGE1_IND[72] <= 8'd18;
    STAGE1_IND[73] <= 8'd146;
    STAGE1_IND[74] <= 8'd82;
    STAGE1_IND[75] <= 8'd210;
    STAGE1_IND[76] <= 8'd50;
    STAGE1_IND[77] <= 8'd178;
    STAGE1_IND[78] <= 8'd114;
    STAGE1_IND[79] <= 8'd242;
    STAGE1_IND[80] <= 8'd10;
    STAGE1_IND[81] <= 8'd138;
    STAGE1_IND[82] <= 8'd74;
    STAGE1_IND[83] <= 8'd202;
    STAGE1_IND[84] <= 8'd42;
    STAGE1_IND[85] <= 8'd170;
    STAGE1_IND[86] <= 8'd106;
    STAGE1_IND[87] <= 8'd234;
    STAGE1_IND[88] <= 8'd26;
    STAGE1_IND[89] <= 8'd154;
    STAGE1_IND[90] <= 8'd90;
    STAGE1_IND[91] <= 8'd218;
    STAGE1_IND[92] <= 8'd58;
    STAGE1_IND[93] <= 8'd186;
    STAGE1_IND[94] <= 8'd122;
    STAGE1_IND[95] <= 8'd250;
    STAGE1_IND[96] <= 8'd6;
    STAGE1_IND[97] <= 8'd134;
    STAGE1_IND[98] <= 8'd70;
    STAGE1_IND[99] <= 8'd198;
    STAGE1_IND[100] <= 8'd38;
    STAGE1_IND[101] <= 8'd166;
    STAGE1_IND[102] <= 8'd102;
    STAGE1_IND[103] <= 8'd230;
    STAGE1_IND[104] <= 8'd22;
    STAGE1_IND[105] <= 8'd150;
    STAGE1_IND[106] <= 8'd86;
    STAGE1_IND[107] <= 8'd214;
    STAGE1_IND[108] <= 8'd54;
    STAGE1_IND[109] <= 8'd182;
    STAGE1_IND[110] <= 8'd118;
    STAGE1_IND[111] <= 8'd246;
    STAGE1_IND[112] <= 8'd14;
    STAGE1_IND[113] <= 8'd142;
    STAGE1_IND[114] <= 8'd78;
    STAGE1_IND[115] <= 8'd206;
    STAGE1_IND[116] <= 8'd46;
    STAGE1_IND[117] <= 8'd174;
    STAGE1_IND[118] <= 8'd110;
    STAGE1_IND[119] <= 8'd238;
    STAGE1_IND[120] <= 8'd30;
    STAGE1_IND[121] <= 8'd158;
    STAGE1_IND[122] <= 8'd94;
    STAGE1_IND[123] <= 8'd222;
    STAGE1_IND[124] <= 8'd62;
    STAGE1_IND[125] <= 8'd190;
    STAGE1_IND[126] <= 8'd126;
    STAGE1_IND[127] <= 8'd254;
    STAGE1_IND[128] <= 8'd1;
    STAGE1_IND[129] <= 8'd129;
    STAGE1_IND[130] <= 8'd65;
    STAGE1_IND[131] <= 8'd193;
    STAGE1_IND[132] <= 8'd33;
    STAGE1_IND[133] <= 8'd161;
    STAGE1_IND[134] <= 8'd97;
    STAGE1_IND[135] <= 8'd225;
    STAGE1_IND[136] <= 8'd17;
    STAGE1_IND[137] <= 8'd145;
    STAGE1_IND[138] <= 8'd81;
    STAGE1_IND[139] <= 8'd209;
    STAGE1_IND[140] <= 8'd49;
    STAGE1_IND[141] <= 8'd177;
    STAGE1_IND[142] <= 8'd113;
    STAGE1_IND[143] <= 8'd241;
    STAGE1_IND[144] <= 8'd9;
    STAGE1_IND[145] <= 8'd137;
    STAGE1_IND[146] <= 8'd73;
    STAGE1_IND[147] <= 8'd201;
    STAGE1_IND[148] <= 8'd41;
    STAGE1_IND[149] <= 8'd169;
    STAGE1_IND[150] <= 8'd105;
    STAGE1_IND[151] <= 8'd233;
    STAGE1_IND[152] <= 8'd25;
    STAGE1_IND[153] <= 8'd153;
    STAGE1_IND[154] <= 8'd89;
    STAGE1_IND[155] <= 8'd217;
    STAGE1_IND[156] <= 8'd57;
    STAGE1_IND[157] <= 8'd185;
    STAGE1_IND[158] <= 8'd121;
    STAGE1_IND[159] <= 8'd249;
    STAGE1_IND[160] <= 8'd5;
    STAGE1_IND[161] <= 8'd133;
    STAGE1_IND[162] <= 8'd69;
    STAGE1_IND[163] <= 8'd197;
    STAGE1_IND[164] <= 8'd37;
    STAGE1_IND[165] <= 8'd165;
    STAGE1_IND[166] <= 8'd101;
    STAGE1_IND[167] <= 8'd229;
    STAGE1_IND[168] <= 8'd21;
    STAGE1_IND[169] <= 8'd149;
    STAGE1_IND[170] <= 8'd85;
    STAGE1_IND[171] <= 8'd213;
    STAGE1_IND[172] <= 8'd53;
    STAGE1_IND[173] <= 8'd181;
    STAGE1_IND[174] <= 8'd117;
    STAGE1_IND[175] <= 8'd245;
    STAGE1_IND[176] <= 8'd13;
    STAGE1_IND[177] <= 8'd141;
    STAGE1_IND[178] <= 8'd77;
    STAGE1_IND[179] <= 8'd205;
    STAGE1_IND[180] <= 8'd45;
    STAGE1_IND[181] <= 8'd173;
    STAGE1_IND[182] <= 8'd109;
    STAGE1_IND[183] <= 8'd237;
    STAGE1_IND[184] <= 8'd29;
    STAGE1_IND[185] <= 8'd157;
    STAGE1_IND[186] <= 8'd93;
    STAGE1_IND[187] <= 8'd221;
    STAGE1_IND[188] <= 8'd61;
    STAGE1_IND[189] <= 8'd189;
    STAGE1_IND[190] <= 8'd125;
    STAGE1_IND[191] <= 8'd253;
    STAGE1_IND[192] <= 8'd3;
    STAGE1_IND[193] <= 8'd131;
    STAGE1_IND[194] <= 8'd67;
    STAGE1_IND[195] <= 8'd195;
    STAGE1_IND[196] <= 8'd35;
    STAGE1_IND[197] <= 8'd163;
    STAGE1_IND[198] <= 8'd99;
    STAGE1_IND[199] <= 8'd227;
    STAGE1_IND[200] <= 8'd19;
    STAGE1_IND[201] <= 8'd147;
    STAGE1_IND[202] <= 8'd83;
    STAGE1_IND[203] <= 8'd211;
    STAGE1_IND[204] <= 8'd51;
    STAGE1_IND[205] <= 8'd179;
    STAGE1_IND[206] <= 8'd115;
    STAGE1_IND[207] <= 8'd243;
    STAGE1_IND[208] <= 8'd11;
    STAGE1_IND[209] <= 8'd139;
    STAGE1_IND[210] <= 8'd75;
    STAGE1_IND[211] <= 8'd203;
    STAGE1_IND[212] <= 8'd43;
    STAGE1_IND[213] <= 8'd171;
    STAGE1_IND[214] <= 8'd107;
    STAGE1_IND[215] <= 8'd235;
    STAGE1_IND[216] <= 8'd27;
    STAGE1_IND[217] <= 8'd155;
    STAGE1_IND[218] <= 8'd91;
    STAGE1_IND[219] <= 8'd219;
    STAGE1_IND[220] <= 8'd59;
    STAGE1_IND[221] <= 8'd187;
    STAGE1_IND[222] <= 8'd123;
    STAGE1_IND[223] <= 8'd251;
    STAGE1_IND[224] <= 8'd7;
    STAGE1_IND[225] <= 8'd135;
    STAGE1_IND[226] <= 8'd71;
    STAGE1_IND[227] <= 8'd199;
    STAGE1_IND[228] <= 8'd39;
    STAGE1_IND[229] <= 8'd167;
    STAGE1_IND[230] <= 8'd103;
    STAGE1_IND[231] <= 8'd231;
    STAGE1_IND[232] <= 8'd23;
    STAGE1_IND[233] <= 8'd151;
    STAGE1_IND[234] <= 8'd87;
    STAGE1_IND[235] <= 8'd215;
    STAGE1_IND[236] <= 8'd55;
    STAGE1_IND[237] <= 8'd183;
    STAGE1_IND[238] <= 8'd119;
    STAGE1_IND[239] <= 8'd247;
    STAGE1_IND[240] <= 8'd15;
    STAGE1_IND[241] <= 8'd143;
    STAGE1_IND[242] <= 8'd79;
    STAGE1_IND[243] <= 8'd207;
    STAGE1_IND[244] <= 8'd47;
    STAGE1_IND[245] <= 8'd175;
    STAGE1_IND[246] <= 8'd111;
    STAGE1_IND[247] <= 8'd239;
    STAGE1_IND[248] <= 8'd31;
    STAGE1_IND[249] <= 8'd159;
    STAGE1_IND[250] <= 8'd95;
    STAGE1_IND[251] <= 8'd223;
    STAGE1_IND[252] <= 8'd63;
    STAGE1_IND[253] <= 8'd191;
    STAGE1_IND[254] <= 8'd127;
    STAGE1_IND[255] <= 8'd255;
end
initial begin
       STAGE2_IND[0] <= 8'd0;
    STAGE2_IND[1] <= 8'd64;
    STAGE2_IND[2] <= 8'd128;
    STAGE2_IND[3] <= 8'd192;
    STAGE2_IND[4] <= 8'd32;
    STAGE2_IND[5] <= 8'd96;
    STAGE2_IND[6] <= 8'd160;
    STAGE2_IND[7] <= 8'd224;
    STAGE2_IND[8] <= 8'd16;
    STAGE2_IND[9] <= 8'd80;
    STAGE2_IND[10] <= 8'd144;
    STAGE2_IND[11] <= 8'd208;
    STAGE2_IND[12] <= 8'd48;
    STAGE2_IND[13] <= 8'd112;
    STAGE2_IND[14] <= 8'd176;
    STAGE2_IND[15] <= 8'd240;
    STAGE2_IND[16] <= 8'd8;
    STAGE2_IND[17] <= 8'd72;
    STAGE2_IND[18] <= 8'd136;
    STAGE2_IND[19] <= 8'd200;
    STAGE2_IND[20] <= 8'd40;
    STAGE2_IND[21] <= 8'd104;
    STAGE2_IND[22] <= 8'd168;
    STAGE2_IND[23] <= 8'd232;
    STAGE2_IND[24] <= 8'd24;
    STAGE2_IND[25] <= 8'd88;
    STAGE2_IND[26] <= 8'd152;
    STAGE2_IND[27] <= 8'd216;
    STAGE2_IND[28] <= 8'd56;
    STAGE2_IND[29] <= 8'd120;
    STAGE2_IND[30] <= 8'd184;
    STAGE2_IND[31] <= 8'd248;
    STAGE2_IND[32] <= 8'd4;
    STAGE2_IND[33] <= 8'd68;
    STAGE2_IND[34] <= 8'd132;
    STAGE2_IND[35] <= 8'd196;
    STAGE2_IND[36] <= 8'd36;
    STAGE2_IND[37] <= 8'd100;
    STAGE2_IND[38] <= 8'd164;
    STAGE2_IND[39] <= 8'd228;
    STAGE2_IND[40] <= 8'd20;
    STAGE2_IND[41] <= 8'd84;
    STAGE2_IND[42] <= 8'd148;
    STAGE2_IND[43] <= 8'd212;
    STAGE2_IND[44] <= 8'd52;
    STAGE2_IND[45] <= 8'd116;
    STAGE2_IND[46] <= 8'd180;
    STAGE2_IND[47] <= 8'd244;
    STAGE2_IND[48] <= 8'd12;
    STAGE2_IND[49] <= 8'd76;
    STAGE2_IND[50] <= 8'd140;
    STAGE2_IND[51] <= 8'd204;
    STAGE2_IND[52] <= 8'd44;
    STAGE2_IND[53] <= 8'd108;
    STAGE2_IND[54] <= 8'd172;
    STAGE2_IND[55] <= 8'd236;
    STAGE2_IND[56] <= 8'd28;
    STAGE2_IND[57] <= 8'd92;
    STAGE2_IND[58] <= 8'd156;
    STAGE2_IND[59] <= 8'd220;
    STAGE2_IND[60] <= 8'd60;
    STAGE2_IND[61] <= 8'd124;
    STAGE2_IND[62] <= 8'd188;
    STAGE2_IND[63] <= 8'd252;
    STAGE2_IND[64] <= 8'd2;
    STAGE2_IND[65] <= 8'd66;
    STAGE2_IND[66] <= 8'd130;
    STAGE2_IND[67] <= 8'd194;
    STAGE2_IND[68] <= 8'd34;
    STAGE2_IND[69] <= 8'd98;
    STAGE2_IND[70] <= 8'd162;
    STAGE2_IND[71] <= 8'd226;
    STAGE2_IND[72] <= 8'd18;
    STAGE2_IND[73] <= 8'd82;
    STAGE2_IND[74] <= 8'd146;
    STAGE2_IND[75] <= 8'd210;
    STAGE2_IND[76] <= 8'd50;
    STAGE2_IND[77] <= 8'd114;
    STAGE2_IND[78] <= 8'd178;
    STAGE2_IND[79] <= 8'd242;
    STAGE2_IND[80] <= 8'd10;
    STAGE2_IND[81] <= 8'd74;
    STAGE2_IND[82] <= 8'd138;
    STAGE2_IND[83] <= 8'd202;
    STAGE2_IND[84] <= 8'd42;
    STAGE2_IND[85] <= 8'd106;
    STAGE2_IND[86] <= 8'd170;
    STAGE2_IND[87] <= 8'd234;
    STAGE2_IND[88] <= 8'd26;
    STAGE2_IND[89] <= 8'd90;
    STAGE2_IND[90] <= 8'd154;
    STAGE2_IND[91] <= 8'd218;
    STAGE2_IND[92] <= 8'd58;
    STAGE2_IND[93] <= 8'd122;
    STAGE2_IND[94] <= 8'd186;
    STAGE2_IND[95] <= 8'd250;
    STAGE2_IND[96] <= 8'd6;
    STAGE2_IND[97] <= 8'd70;
    STAGE2_IND[98] <= 8'd134;
    STAGE2_IND[99] <= 8'd198;
    STAGE2_IND[100] <= 8'd38;
    STAGE2_IND[101] <= 8'd102;
    STAGE2_IND[102] <= 8'd166;
    STAGE2_IND[103] <= 8'd230;
    STAGE2_IND[104] <= 8'd22;
    STAGE2_IND[105] <= 8'd86;
    STAGE2_IND[106] <= 8'd150;
    STAGE2_IND[107] <= 8'd214;
    STAGE2_IND[108] <= 8'd54;
    STAGE2_IND[109] <= 8'd118;
    STAGE2_IND[110] <= 8'd182;
    STAGE2_IND[111] <= 8'd246;
    STAGE2_IND[112] <= 8'd14;
    STAGE2_IND[113] <= 8'd78;
    STAGE2_IND[114] <= 8'd142;
    STAGE2_IND[115] <= 8'd206;
    STAGE2_IND[116] <= 8'd46;
    STAGE2_IND[117] <= 8'd110;
    STAGE2_IND[118] <= 8'd174;
    STAGE2_IND[119] <= 8'd238;
    STAGE2_IND[120] <= 8'd30;
    STAGE2_IND[121] <= 8'd94;
    STAGE2_IND[122] <= 8'd158;
    STAGE2_IND[123] <= 8'd222;
    STAGE2_IND[124] <= 8'd62;
    STAGE2_IND[125] <= 8'd126;
    STAGE2_IND[126] <= 8'd190;
    STAGE2_IND[127] <= 8'd254;
    STAGE2_IND[128] <= 8'd1;
    STAGE2_IND[129] <= 8'd65;
    STAGE2_IND[130] <= 8'd129;
    STAGE2_IND[131] <= 8'd193;
    STAGE2_IND[132] <= 8'd33;
    STAGE2_IND[133] <= 8'd97;
    STAGE2_IND[134] <= 8'd161;
    STAGE2_IND[135] <= 8'd225;
    STAGE2_IND[136] <= 8'd17;
    STAGE2_IND[137] <= 8'd81;
    STAGE2_IND[138] <= 8'd145;
    STAGE2_IND[139] <= 8'd209;
    STAGE2_IND[140] <= 8'd49;
    STAGE2_IND[141] <= 8'd113;
    STAGE2_IND[142] <= 8'd177;
    STAGE2_IND[143] <= 8'd241;
    STAGE2_IND[144] <= 8'd9;
    STAGE2_IND[145] <= 8'd73;
    STAGE2_IND[146] <= 8'd137;
    STAGE2_IND[147] <= 8'd201;
    STAGE2_IND[148] <= 8'd41;
    STAGE2_IND[149] <= 8'd105;
    STAGE2_IND[150] <= 8'd169;
    STAGE2_IND[151] <= 8'd233;
    STAGE2_IND[152] <= 8'd25;
    STAGE2_IND[153] <= 8'd89;
    STAGE2_IND[154] <= 8'd153;
    STAGE2_IND[155] <= 8'd217;
    STAGE2_IND[156] <= 8'd57;
    STAGE2_IND[157] <= 8'd121;
    STAGE2_IND[158] <= 8'd185;
    STAGE2_IND[159] <= 8'd249;
    STAGE2_IND[160] <= 8'd5;
    STAGE2_IND[161] <= 8'd69;
    STAGE2_IND[162] <= 8'd133;
    STAGE2_IND[163] <= 8'd197;
    STAGE2_IND[164] <= 8'd37;
    STAGE2_IND[165] <= 8'd101;
    STAGE2_IND[166] <= 8'd165;
    STAGE2_IND[167] <= 8'd229;
    STAGE2_IND[168] <= 8'd21;
    STAGE2_IND[169] <= 8'd85;
    STAGE2_IND[170] <= 8'd149;
    STAGE2_IND[171] <= 8'd213;
    STAGE2_IND[172] <= 8'd53;
    STAGE2_IND[173] <= 8'd117;
    STAGE2_IND[174] <= 8'd181;
    STAGE2_IND[175] <= 8'd245;
    STAGE2_IND[176] <= 8'd13;
    STAGE2_IND[177] <= 8'd77;
    STAGE2_IND[178] <= 8'd141;
    STAGE2_IND[179] <= 8'd205;
    STAGE2_IND[180] <= 8'd45;
    STAGE2_IND[181] <= 8'd109;
    STAGE2_IND[182] <= 8'd173;
    STAGE2_IND[183] <= 8'd237;
    STAGE2_IND[184] <= 8'd29;
    STAGE2_IND[185] <= 8'd93;
    STAGE2_IND[186] <= 8'd157;
    STAGE2_IND[187] <= 8'd221;
    STAGE2_IND[188] <= 8'd61;
    STAGE2_IND[189] <= 8'd125;
    STAGE2_IND[190] <= 8'd189;
    STAGE2_IND[191] <= 8'd253;
    STAGE2_IND[192] <= 8'd3;
    STAGE2_IND[193] <= 8'd67;
    STAGE2_IND[194] <= 8'd131;
    STAGE2_IND[195] <= 8'd195;
    STAGE2_IND[196] <= 8'd35;
    STAGE2_IND[197] <= 8'd99;
    STAGE2_IND[198] <= 8'd163;
    STAGE2_IND[199] <= 8'd227;
    STAGE2_IND[200] <= 8'd19;
    STAGE2_IND[201] <= 8'd83;
    STAGE2_IND[202] <= 8'd147;
    STAGE2_IND[203] <= 8'd211;
    STAGE2_IND[204] <= 8'd51;
    STAGE2_IND[205] <= 8'd115;
    STAGE2_IND[206] <= 8'd179;
    STAGE2_IND[207] <= 8'd243;
    STAGE2_IND[208] <= 8'd11;
    STAGE2_IND[209] <= 8'd75;
    STAGE2_IND[210] <= 8'd139;
    STAGE2_IND[211] <= 8'd203;
    STAGE2_IND[212] <= 8'd43;
    STAGE2_IND[213] <= 8'd107;
    STAGE2_IND[214] <= 8'd171;
    STAGE2_IND[215] <= 8'd235;
    STAGE2_IND[216] <= 8'd27;
    STAGE2_IND[217] <= 8'd91;
    STAGE2_IND[218] <= 8'd155;
    STAGE2_IND[219] <= 8'd219;
    STAGE2_IND[220] <= 8'd59;
    STAGE2_IND[221] <= 8'd123;
    STAGE2_IND[222] <= 8'd187;
    STAGE2_IND[223] <= 8'd251;
    STAGE2_IND[224] <= 8'd7;
    STAGE2_IND[225] <= 8'd71;
    STAGE2_IND[226] <= 8'd135;
    STAGE2_IND[227] <= 8'd199;
    STAGE2_IND[228] <= 8'd39;
    STAGE2_IND[229] <= 8'd103;
    STAGE2_IND[230] <= 8'd167;
    STAGE2_IND[231] <= 8'd231;
    STAGE2_IND[232] <= 8'd23;
    STAGE2_IND[233] <= 8'd87;
    STAGE2_IND[234] <= 8'd151;
    STAGE2_IND[235] <= 8'd215;
    STAGE2_IND[236] <= 8'd55;
    STAGE2_IND[237] <= 8'd119;
    STAGE2_IND[238] <= 8'd183;
    STAGE2_IND[239] <= 8'd247;
    STAGE2_IND[240] <= 8'd15;
    STAGE2_IND[241] <= 8'd79;
    STAGE2_IND[242] <= 8'd143;
    STAGE2_IND[243] <= 8'd207;
    STAGE2_IND[244] <= 8'd47;
    STAGE2_IND[245] <= 8'd111;
    STAGE2_IND[246] <= 8'd175;
    STAGE2_IND[247] <= 8'd239;
    STAGE2_IND[248] <= 8'd31;
    STAGE2_IND[249] <= 8'd95;
    STAGE2_IND[250] <= 8'd159;
    STAGE2_IND[251] <= 8'd223;
    STAGE2_IND[252] <= 8'd63;
    STAGE2_IND[253] <= 8'd127;
    STAGE2_IND[254] <= 8'd191;
    STAGE2_IND[255] <= 8'd255;
end
initial begin
        STAGE3_IND[0] <= 8'd0;
    STAGE3_IND[1] <= 8'd32;
    STAGE3_IND[2] <= 8'd128;
    STAGE3_IND[3] <= 8'd160;
    STAGE3_IND[4] <= 8'd64;
    STAGE3_IND[5] <= 8'd96;
    STAGE3_IND[6] <= 8'd192;
    STAGE3_IND[7] <= 8'd224;
    STAGE3_IND[8] <= 8'd16;
    STAGE3_IND[9] <= 8'd48;
    STAGE3_IND[10] <= 8'd144;
    STAGE3_IND[11] <= 8'd176;
    STAGE3_IND[12] <= 8'd80;
    STAGE3_IND[13] <= 8'd112;
    STAGE3_IND[14] <= 8'd208;
    STAGE3_IND[15] <= 8'd240;
    STAGE3_IND[16] <= 8'd8;
    STAGE3_IND[17] <= 8'd40;
    STAGE3_IND[18] <= 8'd136;
    STAGE3_IND[19] <= 8'd168;
    STAGE3_IND[20] <= 8'd72;
    STAGE3_IND[21] <= 8'd104;
    STAGE3_IND[22] <= 8'd200;
    STAGE3_IND[23] <= 8'd232;
    STAGE3_IND[24] <= 8'd24;
    STAGE3_IND[25] <= 8'd56;
    STAGE3_IND[26] <= 8'd152;
    STAGE3_IND[27] <= 8'd184;
    STAGE3_IND[28] <= 8'd88;
    STAGE3_IND[29] <= 8'd120;
    STAGE3_IND[30] <= 8'd216;
    STAGE3_IND[31] <= 8'd248;
    STAGE3_IND[32] <= 8'd4;
    STAGE3_IND[33] <= 8'd36;
    STAGE3_IND[34] <= 8'd132;
    STAGE3_IND[35] <= 8'd164;
    STAGE3_IND[36] <= 8'd68;
    STAGE3_IND[37] <= 8'd100;
    STAGE3_IND[38] <= 8'd196;
    STAGE3_IND[39] <= 8'd228;
    STAGE3_IND[40] <= 8'd20;
    STAGE3_IND[41] <= 8'd52;
    STAGE3_IND[42] <= 8'd148;
    STAGE3_IND[43] <= 8'd180;
    STAGE3_IND[44] <= 8'd84;
    STAGE3_IND[45] <= 8'd116;
    STAGE3_IND[46] <= 8'd212;
    STAGE3_IND[47] <= 8'd244;
    STAGE3_IND[48] <= 8'd12;
    STAGE3_IND[49] <= 8'd44;
    STAGE3_IND[50] <= 8'd140;
    STAGE3_IND[51] <= 8'd172;
    STAGE3_IND[52] <= 8'd76;
    STAGE3_IND[53] <= 8'd108;
    STAGE3_IND[54] <= 8'd204;
    STAGE3_IND[55] <= 8'd236;
    STAGE3_IND[56] <= 8'd28;
    STAGE3_IND[57] <= 8'd60;
    STAGE3_IND[58] <= 8'd156;
    STAGE3_IND[59] <= 8'd188;
    STAGE3_IND[60] <= 8'd92;
    STAGE3_IND[61] <= 8'd124;
    STAGE3_IND[62] <= 8'd220;
    STAGE3_IND[63] <= 8'd252;
    STAGE3_IND[64] <= 8'd2;
    STAGE3_IND[65] <= 8'd34;
    STAGE3_IND[66] <= 8'd130;
    STAGE3_IND[67] <= 8'd162;
    STAGE3_IND[68] <= 8'd66;
    STAGE3_IND[69] <= 8'd98;
    STAGE3_IND[70] <= 8'd194;
    STAGE3_IND[71] <= 8'd226;
    STAGE3_IND[72] <= 8'd18;
    STAGE3_IND[73] <= 8'd50;
    STAGE3_IND[74] <= 8'd146;
    STAGE3_IND[75] <= 8'd178;
    STAGE3_IND[76] <= 8'd82;
    STAGE3_IND[77] <= 8'd114;
    STAGE3_IND[78] <= 8'd210;
    STAGE3_IND[79] <= 8'd242;
    STAGE3_IND[80] <= 8'd10;
    STAGE3_IND[81] <= 8'd42;
    STAGE3_IND[82] <= 8'd138;
    STAGE3_IND[83] <= 8'd170;
    STAGE3_IND[84] <= 8'd74;
    STAGE3_IND[85] <= 8'd106;
    STAGE3_IND[86] <= 8'd202;
    STAGE3_IND[87] <= 8'd234;
    STAGE3_IND[88] <= 8'd26;
    STAGE3_IND[89] <= 8'd58;
    STAGE3_IND[90] <= 8'd154;
    STAGE3_IND[91] <= 8'd186;
    STAGE3_IND[92] <= 8'd90;
    STAGE3_IND[93] <= 8'd122;
    STAGE3_IND[94] <= 8'd218;
    STAGE3_IND[95] <= 8'd250;
    STAGE3_IND[96] <= 8'd6;
    STAGE3_IND[97] <= 8'd38;
    STAGE3_IND[98] <= 8'd134;
    STAGE3_IND[99] <= 8'd166;
    STAGE3_IND[100] <= 8'd70;
    STAGE3_IND[101] <= 8'd102;
    STAGE3_IND[102] <= 8'd198;
    STAGE3_IND[103] <= 8'd230;
    STAGE3_IND[104] <= 8'd22;
    STAGE3_IND[105] <= 8'd54;
    STAGE3_IND[106] <= 8'd150;
    STAGE3_IND[107] <= 8'd182;
    STAGE3_IND[108] <= 8'd86;
    STAGE3_IND[109] <= 8'd118;
    STAGE3_IND[110] <= 8'd214;
    STAGE3_IND[111] <= 8'd246;
    STAGE3_IND[112] <= 8'd14;
    STAGE3_IND[113] <= 8'd46;
    STAGE3_IND[114] <= 8'd142;
    STAGE3_IND[115] <= 8'd174;
    STAGE3_IND[116] <= 8'd78;
    STAGE3_IND[117] <= 8'd110;
    STAGE3_IND[118] <= 8'd206;
    STAGE3_IND[119] <= 8'd238;
    STAGE3_IND[120] <= 8'd30;
    STAGE3_IND[121] <= 8'd62;
    STAGE3_IND[122] <= 8'd158;
    STAGE3_IND[123] <= 8'd190;
    STAGE3_IND[124] <= 8'd94;
    STAGE3_IND[125] <= 8'd126;
    STAGE3_IND[126] <= 8'd222;
    STAGE3_IND[127] <= 8'd254;
    STAGE3_IND[128] <= 8'd1;
    STAGE3_IND[129] <= 8'd33;
    STAGE3_IND[130] <= 8'd129;
    STAGE3_IND[131] <= 8'd161;
    STAGE3_IND[132] <= 8'd65;
    STAGE3_IND[133] <= 8'd97;
    STAGE3_IND[134] <= 8'd193;
    STAGE3_IND[135] <= 8'd225;
    STAGE3_IND[136] <= 8'd17;
    STAGE3_IND[137] <= 8'd49;
    STAGE3_IND[138] <= 8'd145;
    STAGE3_IND[139] <= 8'd177;
    STAGE3_IND[140] <= 8'd81;
    STAGE3_IND[141] <= 8'd113;
    STAGE3_IND[142] <= 8'd209;
    STAGE3_IND[143] <= 8'd241;
    STAGE3_IND[144] <= 8'd9;
    STAGE3_IND[145] <= 8'd41;
    STAGE3_IND[146] <= 8'd137;
    STAGE3_IND[147] <= 8'd169;
    STAGE3_IND[148] <= 8'd73;
    STAGE3_IND[149] <= 8'd105;
    STAGE3_IND[150] <= 8'd201;
    STAGE3_IND[151] <= 8'd233;
    STAGE3_IND[152] <= 8'd25;
    STAGE3_IND[153] <= 8'd57;
    STAGE3_IND[154] <= 8'd153;
    STAGE3_IND[155] <= 8'd185;
    STAGE3_IND[156] <= 8'd89;
    STAGE3_IND[157] <= 8'd121;
    STAGE3_IND[158] <= 8'd217;
    STAGE3_IND[159] <= 8'd249;
    STAGE3_IND[160] <= 8'd5;
    STAGE3_IND[161] <= 8'd37;
    STAGE3_IND[162] <= 8'd133;
    STAGE3_IND[163] <= 8'd165;
    STAGE3_IND[164] <= 8'd69;
    STAGE3_IND[165] <= 8'd101;
    STAGE3_IND[166] <= 8'd197;
    STAGE3_IND[167] <= 8'd229;
    STAGE3_IND[168] <= 8'd21;
    STAGE3_IND[169] <= 8'd53;
    STAGE3_IND[170] <= 8'd149;
    STAGE3_IND[171] <= 8'd181;
    STAGE3_IND[172] <= 8'd85;
    STAGE3_IND[173] <= 8'd117;
    STAGE3_IND[174] <= 8'd213;
    STAGE3_IND[175] <= 8'd245;
    STAGE3_IND[176] <= 8'd13;
    STAGE3_IND[177] <= 8'd45;
    STAGE3_IND[178] <= 8'd141;
    STAGE3_IND[179] <= 8'd173;
    STAGE3_IND[180] <= 8'd77;
    STAGE3_IND[181] <= 8'd109;
    STAGE3_IND[182] <= 8'd205;
    STAGE3_IND[183] <= 8'd237;
    STAGE3_IND[184] <= 8'd29;
    STAGE3_IND[185] <= 8'd61;
    STAGE3_IND[186] <= 8'd157;
    STAGE3_IND[187] <= 8'd189;
    STAGE3_IND[188] <= 8'd93;
    STAGE3_IND[189] <= 8'd125;
    STAGE3_IND[190] <= 8'd221;
    STAGE3_IND[191] <= 8'd253;
    STAGE3_IND[192] <= 8'd3;
    STAGE3_IND[193] <= 8'd35;
    STAGE3_IND[194] <= 8'd131;
    STAGE3_IND[195] <= 8'd163;
    STAGE3_IND[196] <= 8'd67;
    STAGE3_IND[197] <= 8'd99;
    STAGE3_IND[198] <= 8'd195;
    STAGE3_IND[199] <= 8'd227;
    STAGE3_IND[200] <= 8'd19;
    STAGE3_IND[201] <= 8'd51;
    STAGE3_IND[202] <= 8'd147;
    STAGE3_IND[203] <= 8'd179;
    STAGE3_IND[204] <= 8'd83;
    STAGE3_IND[205] <= 8'd115;
    STAGE3_IND[206] <= 8'd211;
    STAGE3_IND[207] <= 8'd243;
    STAGE3_IND[208] <= 8'd11;
    STAGE3_IND[209] <= 8'd43;
    STAGE3_IND[210] <= 8'd139;
    STAGE3_IND[211] <= 8'd171;
    STAGE3_IND[212] <= 8'd75;
    STAGE3_IND[213] <= 8'd107;
    STAGE3_IND[214] <= 8'd203;
    STAGE3_IND[215] <= 8'd235;
    STAGE3_IND[216] <= 8'd27;
    STAGE3_IND[217] <= 8'd59;
    STAGE3_IND[218] <= 8'd155;
    STAGE3_IND[219] <= 8'd187;
    STAGE3_IND[220] <= 8'd91;
    STAGE3_IND[221] <= 8'd123;
    STAGE3_IND[222] <= 8'd219;
    STAGE3_IND[223] <= 8'd251;
    STAGE3_IND[224] <= 8'd7;
    STAGE3_IND[225] <= 8'd39;
    STAGE3_IND[226] <= 8'd135;
    STAGE3_IND[227] <= 8'd167;
    STAGE3_IND[228] <= 8'd71;
    STAGE3_IND[229] <= 8'd103;
    STAGE3_IND[230] <= 8'd199;
    STAGE3_IND[231] <= 8'd231;
    STAGE3_IND[232] <= 8'd23;
    STAGE3_IND[233] <= 8'd55;
    STAGE3_IND[234] <= 8'd151;
    STAGE3_IND[235] <= 8'd183;
    STAGE3_IND[236] <= 8'd87;
    STAGE3_IND[237] <= 8'd119;
    STAGE3_IND[238] <= 8'd215;
    STAGE3_IND[239] <= 8'd247;
    STAGE3_IND[240] <= 8'd15;
    STAGE3_IND[241] <= 8'd47;
    STAGE3_IND[242] <= 8'd143;
    STAGE3_IND[243] <= 8'd175;
    STAGE3_IND[244] <= 8'd79;
    STAGE3_IND[245] <= 8'd111;
    STAGE3_IND[246] <= 8'd207;
    STAGE3_IND[247] <= 8'd239;
    STAGE3_IND[248] <= 8'd31;
    STAGE3_IND[249] <= 8'd63;
    STAGE3_IND[250] <= 8'd159;
    STAGE3_IND[251] <= 8'd191;
    STAGE3_IND[252] <= 8'd95;
    STAGE3_IND[253] <= 8'd127;
    STAGE3_IND[254] <= 8'd223;
    STAGE3_IND[255] <= 8'd255;
end
initial begin
    STAGE4_IND[0] <= 8'd0;
    STAGE4_IND[1] <= 8'd16;
    STAGE4_IND[2] <= 8'd128;
    STAGE4_IND[3] <= 8'd144;
    STAGE4_IND[4] <= 8'd64;
    STAGE4_IND[5] <= 8'd80;
    STAGE4_IND[6] <= 8'd192;
    STAGE4_IND[7] <= 8'd208;
    STAGE4_IND[8] <= 8'd32;
    STAGE4_IND[9] <= 8'd48;
    STAGE4_IND[10] <= 8'd160;
    STAGE4_IND[11] <= 8'd176;
    STAGE4_IND[12] <= 8'd96;
    STAGE4_IND[13] <= 8'd112;
    STAGE4_IND[14] <= 8'd224;
    STAGE4_IND[15] <= 8'd240;
    STAGE4_IND[16] <= 8'd8;
    STAGE4_IND[17] <= 8'd24;
    STAGE4_IND[18] <= 8'd136;
    STAGE4_IND[19] <= 8'd152;
    STAGE4_IND[20] <= 8'd72;
    STAGE4_IND[21] <= 8'd88;
    STAGE4_IND[22] <= 8'd200;
    STAGE4_IND[23] <= 8'd216;
    STAGE4_IND[24] <= 8'd40;
    STAGE4_IND[25] <= 8'd56;
    STAGE4_IND[26] <= 8'd168;
    STAGE4_IND[27] <= 8'd184;
    STAGE4_IND[28] <= 8'd104;
    STAGE4_IND[29] <= 8'd120;
    STAGE4_IND[30] <= 8'd232;
    STAGE4_IND[31] <= 8'd248;
    STAGE4_IND[32] <= 8'd4;
    STAGE4_IND[33] <= 8'd20;
    STAGE4_IND[34] <= 8'd132;
    STAGE4_IND[35] <= 8'd148;
    STAGE4_IND[36] <= 8'd68;
    STAGE4_IND[37] <= 8'd84;
    STAGE4_IND[38] <= 8'd196;
    STAGE4_IND[39] <= 8'd212;
    STAGE4_IND[40] <= 8'd36;
    STAGE4_IND[41] <= 8'd52;
    STAGE4_IND[42] <= 8'd164;
    STAGE4_IND[43] <= 8'd180;
    STAGE4_IND[44] <= 8'd100;
    STAGE4_IND[45] <= 8'd116;
    STAGE4_IND[46] <= 8'd228;
    STAGE4_IND[47] <= 8'd244;
    STAGE4_IND[48] <= 8'd12;
    STAGE4_IND[49] <= 8'd28;
    STAGE4_IND[50] <= 8'd140;
    STAGE4_IND[51] <= 8'd156;
    STAGE4_IND[52] <= 8'd76;
    STAGE4_IND[53] <= 8'd92;
    STAGE4_IND[54] <= 8'd204;
    STAGE4_IND[55] <= 8'd220;
    STAGE4_IND[56] <= 8'd44;
    STAGE4_IND[57] <= 8'd60;
    STAGE4_IND[58] <= 8'd172;
    STAGE4_IND[59] <= 8'd188;
    STAGE4_IND[60] <= 8'd108;
    STAGE4_IND[61] <= 8'd124;
    STAGE4_IND[62] <= 8'd236;
    STAGE4_IND[63] <= 8'd252;
    STAGE4_IND[64] <= 8'd2;
    STAGE4_IND[65] <= 8'd18;
    STAGE4_IND[66] <= 8'd130;
    STAGE4_IND[67] <= 8'd146;
    STAGE4_IND[68] <= 8'd66;
    STAGE4_IND[69] <= 8'd82;
    STAGE4_IND[70] <= 8'd194;
    STAGE4_IND[71] <= 8'd210;
    STAGE4_IND[72] <= 8'd34;
    STAGE4_IND[73] <= 8'd50;
    STAGE4_IND[74] <= 8'd162;
    STAGE4_IND[75] <= 8'd178;
    STAGE4_IND[76] <= 8'd98;
    STAGE4_IND[77] <= 8'd114;
    STAGE4_IND[78] <= 8'd226;
    STAGE4_IND[79] <= 8'd242;
    STAGE4_IND[80] <= 8'd10;
    STAGE4_IND[81] <= 8'd26;
    STAGE4_IND[82] <= 8'd138;
    STAGE4_IND[83] <= 8'd154;
    STAGE4_IND[84] <= 8'd74;
    STAGE4_IND[85] <= 8'd90;
    STAGE4_IND[86] <= 8'd202;
    STAGE4_IND[87] <= 8'd218;
    STAGE4_IND[88] <= 8'd42;
    STAGE4_IND[89] <= 8'd58;
    STAGE4_IND[90] <= 8'd170;
    STAGE4_IND[91] <= 8'd186;
    STAGE4_IND[92] <= 8'd106;
    STAGE4_IND[93] <= 8'd122;
    STAGE4_IND[94] <= 8'd234;
    STAGE4_IND[95] <= 8'd250;
    STAGE4_IND[96] <= 8'd6;
    STAGE4_IND[97] <= 8'd22;
    STAGE4_IND[98] <= 8'd134;
    STAGE4_IND[99] <= 8'd150;
    STAGE4_IND[100] <= 8'd70;
    STAGE4_IND[101] <= 8'd86;
    STAGE4_IND[102] <= 8'd198;
    STAGE4_IND[103] <= 8'd214;
    STAGE4_IND[104] <= 8'd38;
    STAGE4_IND[105] <= 8'd54;
    STAGE4_IND[106] <= 8'd166;
    STAGE4_IND[107] <= 8'd182;
    STAGE4_IND[108] <= 8'd102;
    STAGE4_IND[109] <= 8'd118;
    STAGE4_IND[110] <= 8'd230;
    STAGE4_IND[111] <= 8'd246;
    STAGE4_IND[112] <= 8'd14;
    STAGE4_IND[113] <= 8'd30;
    STAGE4_IND[114] <= 8'd142;
    STAGE4_IND[115] <= 8'd158;
    STAGE4_IND[116] <= 8'd78;
    STAGE4_IND[117] <= 8'd94;
    STAGE4_IND[118] <= 8'd206;
    STAGE4_IND[119] <= 8'd222;
    STAGE4_IND[120] <= 8'd46;
    STAGE4_IND[121] <= 8'd62;
    STAGE4_IND[122] <= 8'd174;
    STAGE4_IND[123] <= 8'd190;
    STAGE4_IND[124] <= 8'd110;
    STAGE4_IND[125] <= 8'd126;
    STAGE4_IND[126] <= 8'd238;
    STAGE4_IND[127] <= 8'd254;
    STAGE4_IND[128] <= 8'd1;
    STAGE4_IND[129] <= 8'd17;
    STAGE4_IND[130] <= 8'd129;
    STAGE4_IND[131] <= 8'd145;
    STAGE4_IND[132] <= 8'd65;
    STAGE4_IND[133] <= 8'd81;
    STAGE4_IND[134] <= 8'd193;
    STAGE4_IND[135] <= 8'd209;
    STAGE4_IND[136] <= 8'd33;
    STAGE4_IND[137] <= 8'd49;
    STAGE4_IND[138] <= 8'd161;
    STAGE4_IND[139] <= 8'd177;
    STAGE4_IND[140] <= 8'd97;
    STAGE4_IND[141] <= 8'd113;
    STAGE4_IND[142] <= 8'd225;
    STAGE4_IND[143] <= 8'd241;
    STAGE4_IND[144] <= 8'd9;
    STAGE4_IND[145] <= 8'd25;
    STAGE4_IND[146] <= 8'd137;
    STAGE4_IND[147] <= 8'd153;
    STAGE4_IND[148] <= 8'd73;
    STAGE4_IND[149] <= 8'd89;
    STAGE4_IND[150] <= 8'd201;
    STAGE4_IND[151] <= 8'd217;
    STAGE4_IND[152] <= 8'd41;
    STAGE4_IND[153] <= 8'd57;
    STAGE4_IND[154] <= 8'd169;
    STAGE4_IND[155] <= 8'd185;
    STAGE4_IND[156] <= 8'd105;
    STAGE4_IND[157] <= 8'd121;
    STAGE4_IND[158] <= 8'd233;
    STAGE4_IND[159] <= 8'd249;
    STAGE4_IND[160] <= 8'd5;
    STAGE4_IND[161] <= 8'd21;
    STAGE4_IND[162] <= 8'd133;
    STAGE4_IND[163] <= 8'd149;
    STAGE4_IND[164] <= 8'd69;
    STAGE4_IND[165] <= 8'd85;
    STAGE4_IND[166] <= 8'd197;
    STAGE4_IND[167] <= 8'd213;
    STAGE4_IND[168] <= 8'd37;
    STAGE4_IND[169] <= 8'd53;
    STAGE4_IND[170] <= 8'd165;
    STAGE4_IND[171] <= 8'd181;
    STAGE4_IND[172] <= 8'd101;
    STAGE4_IND[173] <= 8'd117;
    STAGE4_IND[174] <= 8'd229;
    STAGE4_IND[175] <= 8'd245;
    STAGE4_IND[176] <= 8'd13;
    STAGE4_IND[177] <= 8'd29;
    STAGE4_IND[178] <= 8'd141;
    STAGE4_IND[179] <= 8'd157;
    STAGE4_IND[180] <= 8'd77;
    STAGE4_IND[181] <= 8'd93;
    STAGE4_IND[182] <= 8'd205;
    STAGE4_IND[183] <= 8'd221;
    STAGE4_IND[184] <= 8'd45;
    STAGE4_IND[185] <= 8'd61;
    STAGE4_IND[186] <= 8'd173;
    STAGE4_IND[187] <= 8'd189;
    STAGE4_IND[188] <= 8'd109;
    STAGE4_IND[189] <= 8'd125;
    STAGE4_IND[190] <= 8'd237;
    STAGE4_IND[191] <= 8'd253;
    STAGE4_IND[192] <= 8'd3;
    STAGE4_IND[193] <= 8'd19;
    STAGE4_IND[194] <= 8'd131;
    STAGE4_IND[195] <= 8'd147;
    STAGE4_IND[196] <= 8'd67;
    STAGE4_IND[197] <= 8'd83;
    STAGE4_IND[198] <= 8'd195;
    STAGE4_IND[199] <= 8'd211;
    STAGE4_IND[200] <= 8'd35;
    STAGE4_IND[201] <= 8'd51;
    STAGE4_IND[202] <= 8'd163;
    STAGE4_IND[203] <= 8'd179;
    STAGE4_IND[204] <= 8'd99;
    STAGE4_IND[205] <= 8'd115;
    STAGE4_IND[206] <= 8'd227;
    STAGE4_IND[207] <= 8'd243;
    STAGE4_IND[208] <= 8'd11;
    STAGE4_IND[209] <= 8'd27;
    STAGE4_IND[210] <= 8'd139;
    STAGE4_IND[211] <= 8'd155;
    STAGE4_IND[212] <= 8'd75;
    STAGE4_IND[213] <= 8'd91;
    STAGE4_IND[214] <= 8'd203;
    STAGE4_IND[215] <= 8'd219;
    STAGE4_IND[216] <= 8'd43;
    STAGE4_IND[217] <= 8'd59;
    STAGE4_IND[218] <= 8'd171;
    STAGE4_IND[219] <= 8'd187;
    STAGE4_IND[220] <= 8'd107;
    STAGE4_IND[221] <= 8'd123;
    STAGE4_IND[222] <= 8'd235;
    STAGE4_IND[223] <= 8'd251;
    STAGE4_IND[224] <= 8'd7;
    STAGE4_IND[225] <= 8'd23;
    STAGE4_IND[226] <= 8'd135;
    STAGE4_IND[227] <= 8'd151;
    STAGE4_IND[228] <= 8'd71;
    STAGE4_IND[229] <= 8'd87;
    STAGE4_IND[230] <= 8'd199;
    STAGE4_IND[231] <= 8'd215;
    STAGE4_IND[232] <= 8'd39;
    STAGE4_IND[233] <= 8'd55;
    STAGE4_IND[234] <= 8'd167;
    STAGE4_IND[235] <= 8'd183;
    STAGE4_IND[236] <= 8'd103;
    STAGE4_IND[237] <= 8'd119;
    STAGE4_IND[238] <= 8'd231;
    STAGE4_IND[239] <= 8'd247;
    STAGE4_IND[240] <= 8'd15;
    STAGE4_IND[241] <= 8'd31;
    STAGE4_IND[242] <= 8'd143;
    STAGE4_IND[243] <= 8'd159;
    STAGE4_IND[244] <= 8'd79;
    STAGE4_IND[245] <= 8'd95;
    STAGE4_IND[246] <= 8'd207;
    STAGE4_IND[247] <= 8'd223;
    STAGE4_IND[248] <= 8'd47;
    STAGE4_IND[249] <= 8'd63;
    STAGE4_IND[250] <= 8'd175;
    STAGE4_IND[251] <= 8'd191;
    STAGE4_IND[252] <= 8'd111;
    STAGE4_IND[253] <= 8'd127;
    STAGE4_IND[254] <= 8'd239;
    STAGE4_IND[255] <= 8'd255;
end
initial begin
        STAGE5_IND[0] <= 8'd0;
    STAGE5_IND[1] <= 8'd8;
    STAGE5_IND[2] <= 8'd128;
    STAGE5_IND[3] <= 8'd136;
    STAGE5_IND[4] <= 8'd64;
    STAGE5_IND[5] <= 8'd72;
    STAGE5_IND[6] <= 8'd192;
    STAGE5_IND[7] <= 8'd200;
    STAGE5_IND[8] <= 8'd32;
    STAGE5_IND[9] <= 8'd40;
    STAGE5_IND[10] <= 8'd160;
    STAGE5_IND[11] <= 8'd168;
    STAGE5_IND[12] <= 8'd96;
    STAGE5_IND[13] <= 8'd104;
    STAGE5_IND[14] <= 8'd224;
    STAGE5_IND[15] <= 8'd232;
    STAGE5_IND[16] <= 8'd16;
    STAGE5_IND[17] <= 8'd24;
    STAGE5_IND[18] <= 8'd144;
    STAGE5_IND[19] <= 8'd152;
    STAGE5_IND[20] <= 8'd80;
    STAGE5_IND[21] <= 8'd88;
    STAGE5_IND[22] <= 8'd208;
    STAGE5_IND[23] <= 8'd216;
    STAGE5_IND[24] <= 8'd48;
    STAGE5_IND[25] <= 8'd56;
    STAGE5_IND[26] <= 8'd176;
    STAGE5_IND[27] <= 8'd184;
    STAGE5_IND[28] <= 8'd112;
    STAGE5_IND[29] <= 8'd120;
    STAGE5_IND[30] <= 8'd240;
    STAGE5_IND[31] <= 8'd248;
    STAGE5_IND[32] <= 8'd4;
    STAGE5_IND[33] <= 8'd12;
    STAGE5_IND[34] <= 8'd132;
    STAGE5_IND[35] <= 8'd140;
    STAGE5_IND[36] <= 8'd68;
    STAGE5_IND[37] <= 8'd76;
    STAGE5_IND[38] <= 8'd196;
    STAGE5_IND[39] <= 8'd204;
    STAGE5_IND[40] <= 8'd36;
    STAGE5_IND[41] <= 8'd44;
    STAGE5_IND[42] <= 8'd164;
    STAGE5_IND[43] <= 8'd172;
    STAGE5_IND[44] <= 8'd100;
    STAGE5_IND[45] <= 8'd108;
    STAGE5_IND[46] <= 8'd228;
    STAGE5_IND[47] <= 8'd236;
    STAGE5_IND[48] <= 8'd20;
    STAGE5_IND[49] <= 8'd28;
    STAGE5_IND[50] <= 8'd148;
    STAGE5_IND[51] <= 8'd156;
    STAGE5_IND[52] <= 8'd84;
    STAGE5_IND[53] <= 8'd92;
    STAGE5_IND[54] <= 8'd212;
    STAGE5_IND[55] <= 8'd220;
    STAGE5_IND[56] <= 8'd52;
    STAGE5_IND[57] <= 8'd60;
    STAGE5_IND[58] <= 8'd180;
    STAGE5_IND[59] <= 8'd188;
    STAGE5_IND[60] <= 8'd116;
    STAGE5_IND[61] <= 8'd124;
    STAGE5_IND[62] <= 8'd244;
    STAGE5_IND[63] <= 8'd252;
    STAGE5_IND[64] <= 8'd2;
    STAGE5_IND[65] <= 8'd10;
    STAGE5_IND[66] <= 8'd130;
    STAGE5_IND[67] <= 8'd138;
    STAGE5_IND[68] <= 8'd66;
    STAGE5_IND[69] <= 8'd74;
    STAGE5_IND[70] <= 8'd194;
    STAGE5_IND[71] <= 8'd202;
    STAGE5_IND[72] <= 8'd34;
    STAGE5_IND[73] <= 8'd42;
    STAGE5_IND[74] <= 8'd162;
    STAGE5_IND[75] <= 8'd170;
    STAGE5_IND[76] <= 8'd98;
    STAGE5_IND[77] <= 8'd106;
    STAGE5_IND[78] <= 8'd226;
    STAGE5_IND[79] <= 8'd234;
    STAGE5_IND[80] <= 8'd18;
    STAGE5_IND[81] <= 8'd26;
    STAGE5_IND[82] <= 8'd146;
    STAGE5_IND[83] <= 8'd154;
    STAGE5_IND[84] <= 8'd82;
    STAGE5_IND[85] <= 8'd90;
    STAGE5_IND[86] <= 8'd210;
    STAGE5_IND[87] <= 8'd218;
    STAGE5_IND[88] <= 8'd50;
    STAGE5_IND[89] <= 8'd58;
    STAGE5_IND[90] <= 8'd178;
    STAGE5_IND[91] <= 8'd186;
    STAGE5_IND[92] <= 8'd114;
    STAGE5_IND[93] <= 8'd122;
    STAGE5_IND[94] <= 8'd242;
    STAGE5_IND[95] <= 8'd250;
    STAGE5_IND[96] <= 8'd6;
    STAGE5_IND[97] <= 8'd14;
    STAGE5_IND[98] <= 8'd134;
    STAGE5_IND[99] <= 8'd142;
    STAGE5_IND[100] <= 8'd70;
    STAGE5_IND[101] <= 8'd78;
    STAGE5_IND[102] <= 8'd198;
    STAGE5_IND[103] <= 8'd206;
    STAGE5_IND[104] <= 8'd38;
    STAGE5_IND[105] <= 8'd46;
    STAGE5_IND[106] <= 8'd166;
    STAGE5_IND[107] <= 8'd174;
    STAGE5_IND[108] <= 8'd102;
    STAGE5_IND[109] <= 8'd110;
    STAGE5_IND[110] <= 8'd230;
    STAGE5_IND[111] <= 8'd238;
    STAGE5_IND[112] <= 8'd22;
    STAGE5_IND[113] <= 8'd30;
    STAGE5_IND[114] <= 8'd150;
    STAGE5_IND[115] <= 8'd158;
    STAGE5_IND[116] <= 8'd86;
    STAGE5_IND[117] <= 8'd94;
    STAGE5_IND[118] <= 8'd214;
    STAGE5_IND[119] <= 8'd222;
    STAGE5_IND[120] <= 8'd54;
    STAGE5_IND[121] <= 8'd62;
    STAGE5_IND[122] <= 8'd182;
    STAGE5_IND[123] <= 8'd190;
    STAGE5_IND[124] <= 8'd118;
    STAGE5_IND[125] <= 8'd126;
    STAGE5_IND[126] <= 8'd246;
    STAGE5_IND[127] <= 8'd254;
    STAGE5_IND[128] <= 8'd1;
    STAGE5_IND[129] <= 8'd9;
    STAGE5_IND[130] <= 8'd129;
    STAGE5_IND[131] <= 8'd137;
    STAGE5_IND[132] <= 8'd65;
    STAGE5_IND[133] <= 8'd73;
    STAGE5_IND[134] <= 8'd193;
    STAGE5_IND[135] <= 8'd201;
    STAGE5_IND[136] <= 8'd33;
    STAGE5_IND[137] <= 8'd41;
    STAGE5_IND[138] <= 8'd161;
    STAGE5_IND[139] <= 8'd169;
    STAGE5_IND[140] <= 8'd97;
    STAGE5_IND[141] <= 8'd105;
    STAGE5_IND[142] <= 8'd225;
    STAGE5_IND[143] <= 8'd233;
    STAGE5_IND[144] <= 8'd17;
    STAGE5_IND[145] <= 8'd25;
    STAGE5_IND[146] <= 8'd145;
    STAGE5_IND[147] <= 8'd153;
    STAGE5_IND[148] <= 8'd81;
    STAGE5_IND[149] <= 8'd89;
    STAGE5_IND[150] <= 8'd209;
    STAGE5_IND[151] <= 8'd217;
    STAGE5_IND[152] <= 8'd49;
    STAGE5_IND[153] <= 8'd57;
    STAGE5_IND[154] <= 8'd177;
    STAGE5_IND[155] <= 8'd185;
    STAGE5_IND[156] <= 8'd113;
    STAGE5_IND[157] <= 8'd121;
    STAGE5_IND[158] <= 8'd241;
    STAGE5_IND[159] <= 8'd249;
    STAGE5_IND[160] <= 8'd5;
    STAGE5_IND[161] <= 8'd13;
    STAGE5_IND[162] <= 8'd133;
    STAGE5_IND[163] <= 8'd141;
    STAGE5_IND[164] <= 8'd69;
    STAGE5_IND[165] <= 8'd77;
    STAGE5_IND[166] <= 8'd197;
    STAGE5_IND[167] <= 8'd205;
    STAGE5_IND[168] <= 8'd37;
    STAGE5_IND[169] <= 8'd45;
    STAGE5_IND[170] <= 8'd165;
    STAGE5_IND[171] <= 8'd173;
    STAGE5_IND[172] <= 8'd101;
    STAGE5_IND[173] <= 8'd109;
    STAGE5_IND[174] <= 8'd229;
    STAGE5_IND[175] <= 8'd237;
    STAGE5_IND[176] <= 8'd21;
    STAGE5_IND[177] <= 8'd29;
    STAGE5_IND[178] <= 8'd149;
    STAGE5_IND[179] <= 8'd157;
    STAGE5_IND[180] <= 8'd85;
    STAGE5_IND[181] <= 8'd93;
    STAGE5_IND[182] <= 8'd213;
    STAGE5_IND[183] <= 8'd221;
    STAGE5_IND[184] <= 8'd53;
    STAGE5_IND[185] <= 8'd61;
    STAGE5_IND[186] <= 8'd181;
    STAGE5_IND[187] <= 8'd189;
    STAGE5_IND[188] <= 8'd117;
    STAGE5_IND[189] <= 8'd125;
    STAGE5_IND[190] <= 8'd245;
    STAGE5_IND[191] <= 8'd253;
    STAGE5_IND[192] <= 8'd3;
    STAGE5_IND[193] <= 8'd11;
    STAGE5_IND[194] <= 8'd131;
    STAGE5_IND[195] <= 8'd139;
    STAGE5_IND[196] <= 8'd67;
    STAGE5_IND[197] <= 8'd75;
    STAGE5_IND[198] <= 8'd195;
    STAGE5_IND[199] <= 8'd203;
    STAGE5_IND[200] <= 8'd35;
    STAGE5_IND[201] <= 8'd43;
    STAGE5_IND[202] <= 8'd163;
    STAGE5_IND[203] <= 8'd171;
    STAGE5_IND[204] <= 8'd99;
    STAGE5_IND[205] <= 8'd107;
    STAGE5_IND[206] <= 8'd227;
    STAGE5_IND[207] <= 8'd235;
    STAGE5_IND[208] <= 8'd19;
    STAGE5_IND[209] <= 8'd27;
    STAGE5_IND[210] <= 8'd147;
    STAGE5_IND[211] <= 8'd155;
    STAGE5_IND[212] <= 8'd83;
    STAGE5_IND[213] <= 8'd91;
    STAGE5_IND[214] <= 8'd211;
    STAGE5_IND[215] <= 8'd219;
    STAGE5_IND[216] <= 8'd51;
    STAGE5_IND[217] <= 8'd59;
    STAGE5_IND[218] <= 8'd179;
    STAGE5_IND[219] <= 8'd187;
    STAGE5_IND[220] <= 8'd115;
    STAGE5_IND[221] <= 8'd123;
    STAGE5_IND[222] <= 8'd243;
    STAGE5_IND[223] <= 8'd251;
    STAGE5_IND[224] <= 8'd7;
    STAGE5_IND[225] <= 8'd15;
    STAGE5_IND[226] <= 8'd135;
    STAGE5_IND[227] <= 8'd143;
    STAGE5_IND[228] <= 8'd71;
    STAGE5_IND[229] <= 8'd79;
    STAGE5_IND[230] <= 8'd199;
    STAGE5_IND[231] <= 8'd207;
    STAGE5_IND[232] <= 8'd39;
    STAGE5_IND[233] <= 8'd47;
    STAGE5_IND[234] <= 8'd167;
    STAGE5_IND[235] <= 8'd175;
    STAGE5_IND[236] <= 8'd103;
    STAGE5_IND[237] <= 8'd111;
    STAGE5_IND[238] <= 8'd231;
    STAGE5_IND[239] <= 8'd239;
    STAGE5_IND[240] <= 8'd23;
    STAGE5_IND[241] <= 8'd31;
    STAGE5_IND[242] <= 8'd151;
    STAGE5_IND[243] <= 8'd159;
    STAGE5_IND[244] <= 8'd87;
    STAGE5_IND[245] <= 8'd95;
    STAGE5_IND[246] <= 8'd215;
    STAGE5_IND[247] <= 8'd223;
    STAGE5_IND[248] <= 8'd55;
    STAGE5_IND[249] <= 8'd63;
    STAGE5_IND[250] <= 8'd183;
    STAGE5_IND[251] <= 8'd191;
    STAGE5_IND[252] <= 8'd119;
    STAGE5_IND[253] <= 8'd127;
    STAGE5_IND[254] <= 8'd247;
    STAGE5_IND[255] <= 8'd255;
end
initial begin
    STAGE6_IND[0] <= 8'd0;
    STAGE6_IND[1] <= 8'd4;
    STAGE6_IND[2] <= 8'd128;
    STAGE6_IND[3] <= 8'd132;
    STAGE6_IND[4] <= 8'd64;
    STAGE6_IND[5] <= 8'd68;
    STAGE6_IND[6] <= 8'd192;
    STAGE6_IND[7] <= 8'd196;
    STAGE6_IND[8] <= 8'd32;
    STAGE6_IND[9] <= 8'd36;
    STAGE6_IND[10] <= 8'd160;
    STAGE6_IND[11] <= 8'd164;
    STAGE6_IND[12] <= 8'd96;
    STAGE6_IND[13] <= 8'd100;
    STAGE6_IND[14] <= 8'd224;
    STAGE6_IND[15] <= 8'd228;
    STAGE6_IND[16] <= 8'd16;
    STAGE6_IND[17] <= 8'd20;
    STAGE6_IND[18] <= 8'd144;
    STAGE6_IND[19] <= 8'd148;
    STAGE6_IND[20] <= 8'd80;
    STAGE6_IND[21] <= 8'd84;
    STAGE6_IND[22] <= 8'd208;
    STAGE6_IND[23] <= 8'd212;
    STAGE6_IND[24] <= 8'd48;
    STAGE6_IND[25] <= 8'd52;
    STAGE6_IND[26] <= 8'd176;
    STAGE6_IND[27] <= 8'd180;
    STAGE6_IND[28] <= 8'd112;
    STAGE6_IND[29] <= 8'd116;
    STAGE6_IND[30] <= 8'd240;
    STAGE6_IND[31] <= 8'd244;
    STAGE6_IND[32] <= 8'd8;
    STAGE6_IND[33] <= 8'd12;
    STAGE6_IND[34] <= 8'd136;
    STAGE6_IND[35] <= 8'd140;
    STAGE6_IND[36] <= 8'd72;
    STAGE6_IND[37] <= 8'd76;
    STAGE6_IND[38] <= 8'd200;
    STAGE6_IND[39] <= 8'd204;
    STAGE6_IND[40] <= 8'd40;
    STAGE6_IND[41] <= 8'd44;
    STAGE6_IND[42] <= 8'd168;
    STAGE6_IND[43] <= 8'd172;
    STAGE6_IND[44] <= 8'd104;
    STAGE6_IND[45] <= 8'd108;
    STAGE6_IND[46] <= 8'd232;
    STAGE6_IND[47] <= 8'd236;
    STAGE6_IND[48] <= 8'd24;
    STAGE6_IND[49] <= 8'd28;
    STAGE6_IND[50] <= 8'd152;
    STAGE6_IND[51] <= 8'd156;
    STAGE6_IND[52] <= 8'd88;
    STAGE6_IND[53] <= 8'd92;
    STAGE6_IND[54] <= 8'd216;
    STAGE6_IND[55] <= 8'd220;
    STAGE6_IND[56] <= 8'd56;
    STAGE6_IND[57] <= 8'd60;
    STAGE6_IND[58] <= 8'd184;
    STAGE6_IND[59] <= 8'd188;
    STAGE6_IND[60] <= 8'd120;
    STAGE6_IND[61] <= 8'd124;
    STAGE6_IND[62] <= 8'd248;
    STAGE6_IND[63] <= 8'd252;
    STAGE6_IND[64] <= 8'd2;
    STAGE6_IND[65] <= 8'd6;
    STAGE6_IND[66] <= 8'd130;
    STAGE6_IND[67] <= 8'd134;
    STAGE6_IND[68] <= 8'd66;
    STAGE6_IND[69] <= 8'd70;
    STAGE6_IND[70] <= 8'd194;
    STAGE6_IND[71] <= 8'd198;
    STAGE6_IND[72] <= 8'd34;
    STAGE6_IND[73] <= 8'd38;
    STAGE6_IND[74] <= 8'd162;
    STAGE6_IND[75] <= 8'd166;
    STAGE6_IND[76] <= 8'd98;
    STAGE6_IND[77] <= 8'd102;
    STAGE6_IND[78] <= 8'd226;
    STAGE6_IND[79] <= 8'd230;
    STAGE6_IND[80] <= 8'd18;
    STAGE6_IND[81] <= 8'd22;
    STAGE6_IND[82] <= 8'd146;
    STAGE6_IND[83] <= 8'd150;
    STAGE6_IND[84] <= 8'd82;
    STAGE6_IND[85] <= 8'd86;
    STAGE6_IND[86] <= 8'd210;
    STAGE6_IND[87] <= 8'd214;
    STAGE6_IND[88] <= 8'd50;
    STAGE6_IND[89] <= 8'd54;
    STAGE6_IND[90] <= 8'd178;
    STAGE6_IND[91] <= 8'd182;
    STAGE6_IND[92] <= 8'd114;
    STAGE6_IND[93] <= 8'd118;
    STAGE6_IND[94] <= 8'd242;
    STAGE6_IND[95] <= 8'd246;
    STAGE6_IND[96] <= 8'd10;
    STAGE6_IND[97] <= 8'd14;
    STAGE6_IND[98] <= 8'd138;
    STAGE6_IND[99] <= 8'd142;
    STAGE6_IND[100] <= 8'd74;
    STAGE6_IND[101] <= 8'd78;
    STAGE6_IND[102] <= 8'd202;
    STAGE6_IND[103] <= 8'd206;
    STAGE6_IND[104] <= 8'd42;
    STAGE6_IND[105] <= 8'd46;
    STAGE6_IND[106] <= 8'd170;
    STAGE6_IND[107] <= 8'd174;
    STAGE6_IND[108] <= 8'd106;
    STAGE6_IND[109] <= 8'd110;
    STAGE6_IND[110] <= 8'd234;
    STAGE6_IND[111] <= 8'd238;
    STAGE6_IND[112] <= 8'd26;
    STAGE6_IND[113] <= 8'd30;
    STAGE6_IND[114] <= 8'd154;
    STAGE6_IND[115] <= 8'd158;
    STAGE6_IND[116] <= 8'd90;
    STAGE6_IND[117] <= 8'd94;
    STAGE6_IND[118] <= 8'd218;
    STAGE6_IND[119] <= 8'd222;
    STAGE6_IND[120] <= 8'd58;
    STAGE6_IND[121] <= 8'd62;
    STAGE6_IND[122] <= 8'd186;
    STAGE6_IND[123] <= 8'd190;
    STAGE6_IND[124] <= 8'd122;
    STAGE6_IND[125] <= 8'd126;
    STAGE6_IND[126] <= 8'd250;
    STAGE6_IND[127] <= 8'd254;
    STAGE6_IND[128] <= 8'd1;
    STAGE6_IND[129] <= 8'd5;
    STAGE6_IND[130] <= 8'd129;
    STAGE6_IND[131] <= 8'd133;
    STAGE6_IND[132] <= 8'd65;
    STAGE6_IND[133] <= 8'd69;
    STAGE6_IND[134] <= 8'd193;
    STAGE6_IND[135] <= 8'd197;
    STAGE6_IND[136] <= 8'd33;
    STAGE6_IND[137] <= 8'd37;
    STAGE6_IND[138] <= 8'd161;
    STAGE6_IND[139] <= 8'd165;
    STAGE6_IND[140] <= 8'd97;
    STAGE6_IND[141] <= 8'd101;
    STAGE6_IND[142] <= 8'd225;
    STAGE6_IND[143] <= 8'd229;
    STAGE6_IND[144] <= 8'd17;
    STAGE6_IND[145] <= 8'd21;
    STAGE6_IND[146] <= 8'd145;
    STAGE6_IND[147] <= 8'd149;
    STAGE6_IND[148] <= 8'd81;
    STAGE6_IND[149] <= 8'd85;
    STAGE6_IND[150] <= 8'd209;
    STAGE6_IND[151] <= 8'd213;
    STAGE6_IND[152] <= 8'd49;
    STAGE6_IND[153] <= 8'd53;
    STAGE6_IND[154] <= 8'd177;
    STAGE6_IND[155] <= 8'd181;
    STAGE6_IND[156] <= 8'd113;
    STAGE6_IND[157] <= 8'd117;
    STAGE6_IND[158] <= 8'd241;
    STAGE6_IND[159] <= 8'd245;
    STAGE6_IND[160] <= 8'd9;
    STAGE6_IND[161] <= 8'd13;
    STAGE6_IND[162] <= 8'd137;
    STAGE6_IND[163] <= 8'd141;
    STAGE6_IND[164] <= 8'd73;
    STAGE6_IND[165] <= 8'd77;
    STAGE6_IND[166] <= 8'd201;
    STAGE6_IND[167] <= 8'd205;
    STAGE6_IND[168] <= 8'd41;
    STAGE6_IND[169] <= 8'd45;
    STAGE6_IND[170] <= 8'd169;
    STAGE6_IND[171] <= 8'd173;
    STAGE6_IND[172] <= 8'd105;
    STAGE6_IND[173] <= 8'd109;
    STAGE6_IND[174] <= 8'd233;
    STAGE6_IND[175] <= 8'd237;
    STAGE6_IND[176] <= 8'd25;
    STAGE6_IND[177] <= 8'd29;
    STAGE6_IND[178] <= 8'd153;
    STAGE6_IND[179] <= 8'd157;
    STAGE6_IND[180] <= 8'd89;
    STAGE6_IND[181] <= 8'd93;
    STAGE6_IND[182] <= 8'd217;
    STAGE6_IND[183] <= 8'd221;
    STAGE6_IND[184] <= 8'd57;
    STAGE6_IND[185] <= 8'd61;
    STAGE6_IND[186] <= 8'd185;
    STAGE6_IND[187] <= 8'd189;
    STAGE6_IND[188] <= 8'd121;
    STAGE6_IND[189] <= 8'd125;
    STAGE6_IND[190] <= 8'd249;
    STAGE6_IND[191] <= 8'd253;
    STAGE6_IND[192] <= 8'd3;
    STAGE6_IND[193] <= 8'd7;
    STAGE6_IND[194] <= 8'd131;
    STAGE6_IND[195] <= 8'd135;
    STAGE6_IND[196] <= 8'd67;
    STAGE6_IND[197] <= 8'd71;
    STAGE6_IND[198] <= 8'd195;
    STAGE6_IND[199] <= 8'd199;
    STAGE6_IND[200] <= 8'd35;
    STAGE6_IND[201] <= 8'd39;
    STAGE6_IND[202] <= 8'd163;
    STAGE6_IND[203] <= 8'd167;
    STAGE6_IND[204] <= 8'd99;
    STAGE6_IND[205] <= 8'd103;
    STAGE6_IND[206] <= 8'd227;
    STAGE6_IND[207] <= 8'd231;
    STAGE6_IND[208] <= 8'd19;
    STAGE6_IND[209] <= 8'd23;
    STAGE6_IND[210] <= 8'd147;
    STAGE6_IND[211] <= 8'd151;
    STAGE6_IND[212] <= 8'd83;
    STAGE6_IND[213] <= 8'd87;
    STAGE6_IND[214] <= 8'd211;
    STAGE6_IND[215] <= 8'd215;
    STAGE6_IND[216] <= 8'd51;
    STAGE6_IND[217] <= 8'd55;
    STAGE6_IND[218] <= 8'd179;
    STAGE6_IND[219] <= 8'd183;
    STAGE6_IND[220] <= 8'd115;
    STAGE6_IND[221] <= 8'd119;
    STAGE6_IND[222] <= 8'd243;
    STAGE6_IND[223] <= 8'd247;
    STAGE6_IND[224] <= 8'd11;
    STAGE6_IND[225] <= 8'd15;
    STAGE6_IND[226] <= 8'd139;
    STAGE6_IND[227] <= 8'd143;
    STAGE6_IND[228] <= 8'd75;
    STAGE6_IND[229] <= 8'd79;
    STAGE6_IND[230] <= 8'd203;
    STAGE6_IND[231] <= 8'd207;
    STAGE6_IND[232] <= 8'd43;
    STAGE6_IND[233] <= 8'd47;
    STAGE6_IND[234] <= 8'd171;
    STAGE6_IND[235] <= 8'd175;
    STAGE6_IND[236] <= 8'd107;
    STAGE6_IND[237] <= 8'd111;
    STAGE6_IND[238] <= 8'd235;
    STAGE6_IND[239] <= 8'd239;
    STAGE6_IND[240] <= 8'd27;
    STAGE6_IND[241] <= 8'd31;
    STAGE6_IND[242] <= 8'd155;
    STAGE6_IND[243] <= 8'd159;
    STAGE6_IND[244] <= 8'd91;
    STAGE6_IND[245] <= 8'd95;
    STAGE6_IND[246] <= 8'd219;
    STAGE6_IND[247] <= 8'd223;
    STAGE6_IND[248] <= 8'd59;
    STAGE6_IND[249] <= 8'd63;
    STAGE6_IND[250] <= 8'd187;
    STAGE6_IND[251] <= 8'd191;
    STAGE6_IND[252] <= 8'd123;
    STAGE6_IND[253] <= 8'd127;
    STAGE6_IND[254] <= 8'd251;
    STAGE6_IND[255] <= 8'd255;
end
initial begin
      STAGE7_IND[0] <= 8'd0;
    STAGE7_IND[1] <= 8'd2;
    STAGE7_IND[2] <= 8'd128;
    STAGE7_IND[3] <= 8'd130;
    STAGE7_IND[4] <= 8'd64;
    STAGE7_IND[5] <= 8'd66;
    STAGE7_IND[6] <= 8'd192;
    STAGE7_IND[7] <= 8'd194;
    STAGE7_IND[8] <= 8'd32;
    STAGE7_IND[9] <= 8'd34;
    STAGE7_IND[10] <= 8'd160;
    STAGE7_IND[11] <= 8'd162;
    STAGE7_IND[12] <= 8'd96;
    STAGE7_IND[13] <= 8'd98;
    STAGE7_IND[14] <= 8'd224;
    STAGE7_IND[15] <= 8'd226;
    STAGE7_IND[16] <= 8'd16;
    STAGE7_IND[17] <= 8'd18;
    STAGE7_IND[18] <= 8'd144;
    STAGE7_IND[19] <= 8'd146;
    STAGE7_IND[20] <= 8'd80;
    STAGE7_IND[21] <= 8'd82;
    STAGE7_IND[22] <= 8'd208;
    STAGE7_IND[23] <= 8'd210;
    STAGE7_IND[24] <= 8'd48;
    STAGE7_IND[25] <= 8'd50;
    STAGE7_IND[26] <= 8'd176;
    STAGE7_IND[27] <= 8'd178;
    STAGE7_IND[28] <= 8'd112;
    STAGE7_IND[29] <= 8'd114;
    STAGE7_IND[30] <= 8'd240;
    STAGE7_IND[31] <= 8'd242;
    STAGE7_IND[32] <= 8'd8;
    STAGE7_IND[33] <= 8'd10;
    STAGE7_IND[34] <= 8'd136;
    STAGE7_IND[35] <= 8'd138;
    STAGE7_IND[36] <= 8'd72;
    STAGE7_IND[37] <= 8'd74;
    STAGE7_IND[38] <= 8'd200;
    STAGE7_IND[39] <= 8'd202;
    STAGE7_IND[40] <= 8'd40;
    STAGE7_IND[41] <= 8'd42;
    STAGE7_IND[42] <= 8'd168;
    STAGE7_IND[43] <= 8'd170;
    STAGE7_IND[44] <= 8'd104;
    STAGE7_IND[45] <= 8'd106;
    STAGE7_IND[46] <= 8'd232;
    STAGE7_IND[47] <= 8'd234;
    STAGE7_IND[48] <= 8'd24;
    STAGE7_IND[49] <= 8'd26;
    STAGE7_IND[50] <= 8'd152;
    STAGE7_IND[51] <= 8'd154;
    STAGE7_IND[52] <= 8'd88;
    STAGE7_IND[53] <= 8'd90;
    STAGE7_IND[54] <= 8'd216;
    STAGE7_IND[55] <= 8'd218;
    STAGE7_IND[56] <= 8'd56;
    STAGE7_IND[57] <= 8'd58;
    STAGE7_IND[58] <= 8'd184;
    STAGE7_IND[59] <= 8'd186;
    STAGE7_IND[60] <= 8'd120;
    STAGE7_IND[61] <= 8'd122;
    STAGE7_IND[62] <= 8'd248;
    STAGE7_IND[63] <= 8'd250;
    STAGE7_IND[64] <= 8'd4;
    STAGE7_IND[65] <= 8'd6;
    STAGE7_IND[66] <= 8'd132;
    STAGE7_IND[67] <= 8'd134;
    STAGE7_IND[68] <= 8'd68;
    STAGE7_IND[69] <= 8'd70;
    STAGE7_IND[70] <= 8'd196;
    STAGE7_IND[71] <= 8'd198;
    STAGE7_IND[72] <= 8'd36;
    STAGE7_IND[73] <= 8'd38;
    STAGE7_IND[74] <= 8'd164;
    STAGE7_IND[75] <= 8'd166;
    STAGE7_IND[76] <= 8'd100;
    STAGE7_IND[77] <= 8'd102;
    STAGE7_IND[78] <= 8'd228;
    STAGE7_IND[79] <= 8'd230;
    STAGE7_IND[80] <= 8'd20;
    STAGE7_IND[81] <= 8'd22;
    STAGE7_IND[82] <= 8'd148;
    STAGE7_IND[83] <= 8'd150;
    STAGE7_IND[84] <= 8'd84;
    STAGE7_IND[85] <= 8'd86;
    STAGE7_IND[86] <= 8'd212;
    STAGE7_IND[87] <= 8'd214;
    STAGE7_IND[88] <= 8'd52;
    STAGE7_IND[89] <= 8'd54;
    STAGE7_IND[90] <= 8'd180;
    STAGE7_IND[91] <= 8'd182;
    STAGE7_IND[92] <= 8'd116;
    STAGE7_IND[93] <= 8'd118;
    STAGE7_IND[94] <= 8'd244;
    STAGE7_IND[95] <= 8'd246;
    STAGE7_IND[96] <= 8'd12;
    STAGE7_IND[97] <= 8'd14;
    STAGE7_IND[98] <= 8'd140;
    STAGE7_IND[99] <= 8'd142;
    STAGE7_IND[100] <= 8'd76;
    STAGE7_IND[101] <= 8'd78;
    STAGE7_IND[102] <= 8'd204;
    STAGE7_IND[103] <= 8'd206;
    STAGE7_IND[104] <= 8'd44;
    STAGE7_IND[105] <= 8'd46;
    STAGE7_IND[106] <= 8'd172;
    STAGE7_IND[107] <= 8'd174;
    STAGE7_IND[108] <= 8'd108;
    STAGE7_IND[109] <= 8'd110;
    STAGE7_IND[110] <= 8'd236;
    STAGE7_IND[111] <= 8'd238;
    STAGE7_IND[112] <= 8'd28;
    STAGE7_IND[113] <= 8'd30;
    STAGE7_IND[114] <= 8'd156;
    STAGE7_IND[115] <= 8'd158;
    STAGE7_IND[116] <= 8'd92;
    STAGE7_IND[117] <= 8'd94;
    STAGE7_IND[118] <= 8'd220;
    STAGE7_IND[119] <= 8'd222;
    STAGE7_IND[120] <= 8'd60;
    STAGE7_IND[121] <= 8'd62;
    STAGE7_IND[122] <= 8'd188;
    STAGE7_IND[123] <= 8'd190;
    STAGE7_IND[124] <= 8'd124;
    STAGE7_IND[125] <= 8'd126;
    STAGE7_IND[126] <= 8'd252;
    STAGE7_IND[127] <= 8'd254;
    STAGE7_IND[128] <= 8'd1;
    STAGE7_IND[129] <= 8'd3;
    STAGE7_IND[130] <= 8'd129;
    STAGE7_IND[131] <= 8'd131;
    STAGE7_IND[132] <= 8'd65;
    STAGE7_IND[133] <= 8'd67;
    STAGE7_IND[134] <= 8'd193;
    STAGE7_IND[135] <= 8'd195;
    STAGE7_IND[136] <= 8'd33;
    STAGE7_IND[137] <= 8'd35;
    STAGE7_IND[138] <= 8'd161;
    STAGE7_IND[139] <= 8'd163;
    STAGE7_IND[140] <= 8'd97;
    STAGE7_IND[141] <= 8'd99;
    STAGE7_IND[142] <= 8'd225;
    STAGE7_IND[143] <= 8'd227;
    STAGE7_IND[144] <= 8'd17;
    STAGE7_IND[145] <= 8'd19;
    STAGE7_IND[146] <= 8'd145;
    STAGE7_IND[147] <= 8'd147;
    STAGE7_IND[148] <= 8'd81;
    STAGE7_IND[149] <= 8'd83;
    STAGE7_IND[150] <= 8'd209;
    STAGE7_IND[151] <= 8'd211;
    STAGE7_IND[152] <= 8'd49;
    STAGE7_IND[153] <= 8'd51;
    STAGE7_IND[154] <= 8'd177;
    STAGE7_IND[155] <= 8'd179;
    STAGE7_IND[156] <= 8'd113;
    STAGE7_IND[157] <= 8'd115;
    STAGE7_IND[158] <= 8'd241;
    STAGE7_IND[159] <= 8'd243;
    STAGE7_IND[160] <= 8'd9;
    STAGE7_IND[161] <= 8'd11;
    STAGE7_IND[162] <= 8'd137;
    STAGE7_IND[163] <= 8'd139;
    STAGE7_IND[164] <= 8'd73;
    STAGE7_IND[165] <= 8'd75;
    STAGE7_IND[166] <= 8'd201;
    STAGE7_IND[167] <= 8'd203;
    STAGE7_IND[168] <= 8'd41;
    STAGE7_IND[169] <= 8'd43;
    STAGE7_IND[170] <= 8'd169;
    STAGE7_IND[171] <= 8'd171;
    STAGE7_IND[172] <= 8'd105;
    STAGE7_IND[173] <= 8'd107;
    STAGE7_IND[174] <= 8'd233;
    STAGE7_IND[175] <= 8'd235;
    STAGE7_IND[176] <= 8'd25;
    STAGE7_IND[177] <= 8'd27;
    STAGE7_IND[178] <= 8'd153;
    STAGE7_IND[179] <= 8'd155;
    STAGE7_IND[180] <= 8'd89;
    STAGE7_IND[181] <= 8'd91;
    STAGE7_IND[182] <= 8'd217;
    STAGE7_IND[183] <= 8'd219;
    STAGE7_IND[184] <= 8'd57;
    STAGE7_IND[185] <= 8'd59;
    STAGE7_IND[186] <= 8'd185;
    STAGE7_IND[187] <= 8'd187;
    STAGE7_IND[188] <= 8'd121;
    STAGE7_IND[189] <= 8'd123;
    STAGE7_IND[190] <= 8'd249;
    STAGE7_IND[191] <= 8'd251;
    STAGE7_IND[192] <= 8'd5;
    STAGE7_IND[193] <= 8'd7;
    STAGE7_IND[194] <= 8'd133;
    STAGE7_IND[195] <= 8'd135;
    STAGE7_IND[196] <= 8'd69;
    STAGE7_IND[197] <= 8'd71;
    STAGE7_IND[198] <= 8'd197;
    STAGE7_IND[199] <= 8'd199;
    STAGE7_IND[200] <= 8'd37;
    STAGE7_IND[201] <= 8'd39;
    STAGE7_IND[202] <= 8'd165;
    STAGE7_IND[203] <= 8'd167;
    STAGE7_IND[204] <= 8'd101;
    STAGE7_IND[205] <= 8'd103;
    STAGE7_IND[206] <= 8'd229;
    STAGE7_IND[207] <= 8'd231;
    STAGE7_IND[208] <= 8'd21;
    STAGE7_IND[209] <= 8'd23;
    STAGE7_IND[210] <= 8'd149;
    STAGE7_IND[211] <= 8'd151;
    STAGE7_IND[212] <= 8'd85;
    STAGE7_IND[213] <= 8'd87;
    STAGE7_IND[214] <= 8'd213;
    STAGE7_IND[215] <= 8'd215;
    STAGE7_IND[216] <= 8'd53;
    STAGE7_IND[217] <= 8'd55;
    STAGE7_IND[218] <= 8'd181;
    STAGE7_IND[219] <= 8'd183;
    STAGE7_IND[220] <= 8'd117;
    STAGE7_IND[221] <= 8'd119;
    STAGE7_IND[222] <= 8'd245;
    STAGE7_IND[223] <= 8'd247;
    STAGE7_IND[224] <= 8'd13;
    STAGE7_IND[225] <= 8'd15;
    STAGE7_IND[226] <= 8'd141;
    STAGE7_IND[227] <= 8'd143;
    STAGE7_IND[228] <= 8'd77;
    STAGE7_IND[229] <= 8'd79;
    STAGE7_IND[230] <= 8'd205;
    STAGE7_IND[231] <= 8'd207;
    STAGE7_IND[232] <= 8'd45;
    STAGE7_IND[233] <= 8'd47;
    STAGE7_IND[234] <= 8'd173;
    STAGE7_IND[235] <= 8'd175;
    STAGE7_IND[236] <= 8'd109;
    STAGE7_IND[237] <= 8'd111;
    STAGE7_IND[238] <= 8'd237;
    STAGE7_IND[239] <= 8'd239;
    STAGE7_IND[240] <= 8'd29;
    STAGE7_IND[241] <= 8'd31;
    STAGE7_IND[242] <= 8'd157;
    STAGE7_IND[243] <= 8'd159;
    STAGE7_IND[244] <= 8'd93;
    STAGE7_IND[245] <= 8'd95;
    STAGE7_IND[246] <= 8'd221;
    STAGE7_IND[247] <= 8'd223;
    STAGE7_IND[248] <= 8'd61;
    STAGE7_IND[249] <= 8'd63;
    STAGE7_IND[250] <= 8'd189;
    STAGE7_IND[251] <= 8'd191;
    STAGE7_IND[252] <= 8'd125;
    STAGE7_IND[253] <= 8'd127;
    STAGE7_IND[254] <= 8'd253;
    STAGE7_IND[255] <= 8'd255;
end
initial begin
    STAGE8_IND[0] <= 8'd0;
    STAGE8_IND[1] <= 8'd1;
    STAGE8_IND[2] <= 8'd128;
    STAGE8_IND[3] <= 8'd129;
    STAGE8_IND[4] <= 8'd64;
    STAGE8_IND[5] <= 8'd65;
    STAGE8_IND[6] <= 8'd192;
    STAGE8_IND[7] <= 8'd193;
    STAGE8_IND[8] <= 8'd32;
    STAGE8_IND[9] <= 8'd33;
    STAGE8_IND[10] <= 8'd160;
    STAGE8_IND[11] <= 8'd161;
    STAGE8_IND[12] <= 8'd96;
    STAGE8_IND[13] <= 8'd97;
    STAGE8_IND[14] <= 8'd224;
    STAGE8_IND[15] <= 8'd225;
    STAGE8_IND[16] <= 8'd16;
    STAGE8_IND[17] <= 8'd17;
    STAGE8_IND[18] <= 8'd144;
    STAGE8_IND[19] <= 8'd145;
    STAGE8_IND[20] <= 8'd80;
    STAGE8_IND[21] <= 8'd81;
    STAGE8_IND[22] <= 8'd208;
    STAGE8_IND[23] <= 8'd209;
    STAGE8_IND[24] <= 8'd48;
    STAGE8_IND[25] <= 8'd49;
    STAGE8_IND[26] <= 8'd176;
    STAGE8_IND[27] <= 8'd177;
    STAGE8_IND[28] <= 8'd112;
    STAGE8_IND[29] <= 8'd113;
    STAGE8_IND[30] <= 8'd240;
    STAGE8_IND[31] <= 8'd241;
    STAGE8_IND[32] <= 8'd8;
    STAGE8_IND[33] <= 8'd9;
    STAGE8_IND[34] <= 8'd136;
    STAGE8_IND[35] <= 8'd137;
    STAGE8_IND[36] <= 8'd72;
    STAGE8_IND[37] <= 8'd73;
    STAGE8_IND[38] <= 8'd200;
    STAGE8_IND[39] <= 8'd201;
    STAGE8_IND[40] <= 8'd40;
    STAGE8_IND[41] <= 8'd41;
    STAGE8_IND[42] <= 8'd168;
    STAGE8_IND[43] <= 8'd169;
    STAGE8_IND[44] <= 8'd104;
    STAGE8_IND[45] <= 8'd105;
    STAGE8_IND[46] <= 8'd232;
    STAGE8_IND[47] <= 8'd233;
    STAGE8_IND[48] <= 8'd24;
    STAGE8_IND[49] <= 8'd25;
    STAGE8_IND[50] <= 8'd152;
    STAGE8_IND[51] <= 8'd153;
    STAGE8_IND[52] <= 8'd88;
    STAGE8_IND[53] <= 8'd89;
    STAGE8_IND[54] <= 8'd216;
    STAGE8_IND[55] <= 8'd217;
    STAGE8_IND[56] <= 8'd56;
    STAGE8_IND[57] <= 8'd57;
    STAGE8_IND[58] <= 8'd184;
    STAGE8_IND[59] <= 8'd185;
    STAGE8_IND[60] <= 8'd120;
    STAGE8_IND[61] <= 8'd121;
    STAGE8_IND[62] <= 8'd248;
    STAGE8_IND[63] <= 8'd249;
    STAGE8_IND[64] <= 8'd4;
    STAGE8_IND[65] <= 8'd5;
    STAGE8_IND[66] <= 8'd132;
    STAGE8_IND[67] <= 8'd133;
    STAGE8_IND[68] <= 8'd68;
    STAGE8_IND[69] <= 8'd69;
    STAGE8_IND[70] <= 8'd196;
    STAGE8_IND[71] <= 8'd197;
    STAGE8_IND[72] <= 8'd36;
    STAGE8_IND[73] <= 8'd37;
    STAGE8_IND[74] <= 8'd164;
    STAGE8_IND[75] <= 8'd165;
    STAGE8_IND[76] <= 8'd100;
    STAGE8_IND[77] <= 8'd101;
    STAGE8_IND[78] <= 8'd228;
    STAGE8_IND[79] <= 8'd229;
    STAGE8_IND[80] <= 8'd20;
    STAGE8_IND[81] <= 8'd21;
    STAGE8_IND[82] <= 8'd148;
    STAGE8_IND[83] <= 8'd149;
    STAGE8_IND[84] <= 8'd84;
    STAGE8_IND[85] <= 8'd85;
    STAGE8_IND[86] <= 8'd212;
    STAGE8_IND[87] <= 8'd213;
    STAGE8_IND[88] <= 8'd52;
    STAGE8_IND[89] <= 8'd53;
    STAGE8_IND[90] <= 8'd180;
    STAGE8_IND[91] <= 8'd181;
    STAGE8_IND[92] <= 8'd116;
    STAGE8_IND[93] <= 8'd117;
    STAGE8_IND[94] <= 8'd244;
    STAGE8_IND[95] <= 8'd245;
    STAGE8_IND[96] <= 8'd12;
    STAGE8_IND[97] <= 8'd13;
    STAGE8_IND[98] <= 8'd140;
    STAGE8_IND[99] <= 8'd141;
    STAGE8_IND[100] <= 8'd76;
    STAGE8_IND[101] <= 8'd77;
    STAGE8_IND[102] <= 8'd204;
    STAGE8_IND[103] <= 8'd205;
    STAGE8_IND[104] <= 8'd44;
    STAGE8_IND[105] <= 8'd45;
    STAGE8_IND[106] <= 8'd172;
    STAGE8_IND[107] <= 8'd173;
    STAGE8_IND[108] <= 8'd108;
    STAGE8_IND[109] <= 8'd109;
    STAGE8_IND[110] <= 8'd236;
    STAGE8_IND[111] <= 8'd237;
    STAGE8_IND[112] <= 8'd28;
    STAGE8_IND[113] <= 8'd29;
    STAGE8_IND[114] <= 8'd156;
    STAGE8_IND[115] <= 8'd157;
    STAGE8_IND[116] <= 8'd92;
    STAGE8_IND[117] <= 8'd93;
    STAGE8_IND[118] <= 8'd220;
    STAGE8_IND[119] <= 8'd221;
    STAGE8_IND[120] <= 8'd60;
    STAGE8_IND[121] <= 8'd61;
    STAGE8_IND[122] <= 8'd188;
    STAGE8_IND[123] <= 8'd189;
    STAGE8_IND[124] <= 8'd124;
    STAGE8_IND[125] <= 8'd125;
    STAGE8_IND[126] <= 8'd252;
    STAGE8_IND[127] <= 8'd253;
    STAGE8_IND[128] <= 8'd2;
    STAGE8_IND[129] <= 8'd3;
    STAGE8_IND[130] <= 8'd130;
    STAGE8_IND[131] <= 8'd131;
    STAGE8_IND[132] <= 8'd66;
    STAGE8_IND[133] <= 8'd67;
    STAGE8_IND[134] <= 8'd194;
    STAGE8_IND[135] <= 8'd195;
    STAGE8_IND[136] <= 8'd34;
    STAGE8_IND[137] <= 8'd35;
    STAGE8_IND[138] <= 8'd162;
    STAGE8_IND[139] <= 8'd163;
    STAGE8_IND[140] <= 8'd98;
    STAGE8_IND[141] <= 8'd99;
    STAGE8_IND[142] <= 8'd226;
    STAGE8_IND[143] <= 8'd227;
    STAGE8_IND[144] <= 8'd18;
    STAGE8_IND[145] <= 8'd19;
    STAGE8_IND[146] <= 8'd146;
    STAGE8_IND[147] <= 8'd147;
    STAGE8_IND[148] <= 8'd82;
    STAGE8_IND[149] <= 8'd83;
    STAGE8_IND[150] <= 8'd210;
    STAGE8_IND[151] <= 8'd211;
    STAGE8_IND[152] <= 8'd50;
    STAGE8_IND[153] <= 8'd51;
    STAGE8_IND[154] <= 8'd178;
    STAGE8_IND[155] <= 8'd179;
    STAGE8_IND[156] <= 8'd114;
    STAGE8_IND[157] <= 8'd115;
    STAGE8_IND[158] <= 8'd242;
    STAGE8_IND[159] <= 8'd243;
    STAGE8_IND[160] <= 8'd10;
    STAGE8_IND[161] <= 8'd11;
    STAGE8_IND[162] <= 8'd138;
    STAGE8_IND[163] <= 8'd139;
    STAGE8_IND[164] <= 8'd74;
    STAGE8_IND[165] <= 8'd75;
    STAGE8_IND[166] <= 8'd202;
    STAGE8_IND[167] <= 8'd203;
    STAGE8_IND[168] <= 8'd42;
    STAGE8_IND[169] <= 8'd43;
    STAGE8_IND[170] <= 8'd170;
    STAGE8_IND[171] <= 8'd171;
    STAGE8_IND[172] <= 8'd106;
    STAGE8_IND[173] <= 8'd107;
    STAGE8_IND[174] <= 8'd234;
    STAGE8_IND[175] <= 8'd235;
    STAGE8_IND[176] <= 8'd26;
    STAGE8_IND[177] <= 8'd27;
    STAGE8_IND[178] <= 8'd154;
    STAGE8_IND[179] <= 8'd155;
    STAGE8_IND[180] <= 8'd90;
    STAGE8_IND[181] <= 8'd91;
    STAGE8_IND[182] <= 8'd218;
    STAGE8_IND[183] <= 8'd219;
    STAGE8_IND[184] <= 8'd58;
    STAGE8_IND[185] <= 8'd59;
    STAGE8_IND[186] <= 8'd186;
    STAGE8_IND[187] <= 8'd187;
    STAGE8_IND[188] <= 8'd122;
    STAGE8_IND[189] <= 8'd123;
    STAGE8_IND[190] <= 8'd250;
    STAGE8_IND[191] <= 8'd251;
    STAGE8_IND[192] <= 8'd6;
    STAGE8_IND[193] <= 8'd7;
    STAGE8_IND[194] <= 8'd134;
    STAGE8_IND[195] <= 8'd135;
    STAGE8_IND[196] <= 8'd70;
    STAGE8_IND[197] <= 8'd71;
    STAGE8_IND[198] <= 8'd198;
    STAGE8_IND[199] <= 8'd199;
    STAGE8_IND[200] <= 8'd38;
    STAGE8_IND[201] <= 8'd39;
    STAGE8_IND[202] <= 8'd166;
    STAGE8_IND[203] <= 8'd167;
    STAGE8_IND[204] <= 8'd102;
    STAGE8_IND[205] <= 8'd103;
    STAGE8_IND[206] <= 8'd230;
    STAGE8_IND[207] <= 8'd231;
    STAGE8_IND[208] <= 8'd22;
    STAGE8_IND[209] <= 8'd23;
    STAGE8_IND[210] <= 8'd150;
    STAGE8_IND[211] <= 8'd151;
    STAGE8_IND[212] <= 8'd86;
    STAGE8_IND[213] <= 8'd87;
    STAGE8_IND[214] <= 8'd214;
    STAGE8_IND[215] <= 8'd215;
    STAGE8_IND[216] <= 8'd54;
    STAGE8_IND[217] <= 8'd55;
    STAGE8_IND[218] <= 8'd182;
    STAGE8_IND[219] <= 8'd183;
    STAGE8_IND[220] <= 8'd118;
    STAGE8_IND[221] <= 8'd119;
    STAGE8_IND[222] <= 8'd246;
    STAGE8_IND[223] <= 8'd247;
    STAGE8_IND[224] <= 8'd14;
    STAGE8_IND[225] <= 8'd15;
    STAGE8_IND[226] <= 8'd142;
    STAGE8_IND[227] <= 8'd143;
    STAGE8_IND[228] <= 8'd78;
    STAGE8_IND[229] <= 8'd79;
    STAGE8_IND[230] <= 8'd206;
    STAGE8_IND[231] <= 8'd207;
    STAGE8_IND[232] <= 8'd46;
    STAGE8_IND[233] <= 8'd47;
    STAGE8_IND[234] <= 8'd174;
    STAGE8_IND[235] <= 8'd175;
    STAGE8_IND[236] <= 8'd110;
    STAGE8_IND[237] <= 8'd111;
    STAGE8_IND[238] <= 8'd238;
    STAGE8_IND[239] <= 8'd239;
    STAGE8_IND[240] <= 8'd30;
    STAGE8_IND[241] <= 8'd31;
    STAGE8_IND[242] <= 8'd158;
    STAGE8_IND[243] <= 8'd159;
    STAGE8_IND[244] <= 8'd94;
    STAGE8_IND[245] <= 8'd95;
    STAGE8_IND[246] <= 8'd222;
    STAGE8_IND[247] <= 8'd223;
    STAGE8_IND[248] <= 8'd62;
    STAGE8_IND[249] <= 8'd63;
    STAGE8_IND[250] <= 8'd190;
    STAGE8_IND[251] <= 8'd191;
    STAGE8_IND[252] <= 8'd126;
    STAGE8_IND[253] <= 8'd127;
    STAGE8_IND[254] <= 8'd254;
    STAGE8_IND[255] <= 8'd255;
end

initial begin
    BITFLIP_IND[0] <= 8'd0;
    BITFLIP_IND[1] <= 8'd1;
    BITFLIP_IND[2] <= 8'd2;
    BITFLIP_IND[3] <= 8'd3;
    BITFLIP_IND[4] <= 8'd4;
    BITFLIP_IND[5] <= 8'd5;
    BITFLIP_IND[6] <= 8'd6;
    BITFLIP_IND[7] <= 8'd7;
    BITFLIP_IND[8] <= 8'd8;
    BITFLIP_IND[9] <= 8'd9;
    BITFLIP_IND[10] <= 8'd10;
    BITFLIP_IND[11] <= 8'd11;
    BITFLIP_IND[12] <= 8'd12;
    BITFLIP_IND[13] <= 8'd13;
    BITFLIP_IND[14] <= 8'd14;
    BITFLIP_IND[15] <= 8'd15;
    BITFLIP_IND[16] <= 8'd16;
    BITFLIP_IND[17] <= 8'd17;
    BITFLIP_IND[18] <= 8'd18;
    BITFLIP_IND[19] <= 8'd19;
    BITFLIP_IND[20] <= 8'd20;
    BITFLIP_IND[21] <= 8'd21;
    BITFLIP_IND[22] <= 8'd22;
    BITFLIP_IND[23] <= 8'd23;
    BITFLIP_IND[24] <= 8'd24;
    BITFLIP_IND[25] <= 8'd25;
    BITFLIP_IND[26] <= 8'd26;
    BITFLIP_IND[27] <= 8'd27;
    BITFLIP_IND[28] <= 8'd28;
    BITFLIP_IND[29] <= 8'd29;
    BITFLIP_IND[30] <= 8'd30;
    BITFLIP_IND[31] <= 8'd31;
    BITFLIP_IND[32] <= 8'd32;
    BITFLIP_IND[33] <= 8'd33;
    BITFLIP_IND[34] <= 8'd34;
    BITFLIP_IND[35] <= 8'd35;
    BITFLIP_IND[36] <= 8'd36;
    BITFLIP_IND[37] <= 8'd37;
    BITFLIP_IND[38] <= 8'd38;
    BITFLIP_IND[39] <= 8'd39;
    BITFLIP_IND[40] <= 8'd40;
    BITFLIP_IND[41] <= 8'd41;
    BITFLIP_IND[42] <= 8'd42;
    BITFLIP_IND[43] <= 8'd43;
    BITFLIP_IND[44] <= 8'd44;
    BITFLIP_IND[45] <= 8'd45;
    BITFLIP_IND[46] <= 8'd46;
    BITFLIP_IND[47] <= 8'd47;
    BITFLIP_IND[48] <= 8'd48;
    BITFLIP_IND[49] <= 8'd49;
    BITFLIP_IND[50] <= 8'd50;
    BITFLIP_IND[51] <= 8'd51;
    BITFLIP_IND[52] <= 8'd52;
    BITFLIP_IND[53] <= 8'd53;
    BITFLIP_IND[54] <= 8'd54;
    BITFLIP_IND[55] <= 8'd55;
    BITFLIP_IND[56] <= 8'd56;
    BITFLIP_IND[57] <= 8'd57;
    BITFLIP_IND[58] <= 8'd58;
    BITFLIP_IND[59] <= 8'd59;
    BITFLIP_IND[60] <= 8'd60;
    BITFLIP_IND[61] <= 8'd61;
    BITFLIP_IND[62] <= 8'd62;
    BITFLIP_IND[63] <= 8'd63;
    BITFLIP_IND[64] <= 8'd64;
    BITFLIP_IND[65] <= 8'd65;
    BITFLIP_IND[66] <= 8'd66;
    BITFLIP_IND[67] <= 8'd67;
    BITFLIP_IND[68] <= 8'd68;
    BITFLIP_IND[69] <= 8'd69;
    BITFLIP_IND[70] <= 8'd70;
    BITFLIP_IND[71] <= 8'd71;
    BITFLIP_IND[72] <= 8'd72;
    BITFLIP_IND[73] <= 8'd73;
    BITFLIP_IND[74] <= 8'd74;
    BITFLIP_IND[75] <= 8'd75;
    BITFLIP_IND[76] <= 8'd76;
    BITFLIP_IND[77] <= 8'd77;
    BITFLIP_IND[78] <= 8'd78;
    BITFLIP_IND[79] <= 8'd79;
    BITFLIP_IND[80] <= 8'd80;
    BITFLIP_IND[81] <= 8'd81;
    BITFLIP_IND[82] <= 8'd82;
    BITFLIP_IND[83] <= 8'd83;
    BITFLIP_IND[84] <= 8'd84;
    BITFLIP_IND[85] <= 8'd85;
    BITFLIP_IND[86] <= 8'd86;
    BITFLIP_IND[87] <= 8'd87;
    BITFLIP_IND[88] <= 8'd88;
    BITFLIP_IND[89] <= 8'd89;
    BITFLIP_IND[90] <= 8'd90;
    BITFLIP_IND[91] <= 8'd91;
    BITFLIP_IND[92] <= 8'd92;
    BITFLIP_IND[93] <= 8'd93;
    BITFLIP_IND[94] <= 8'd94;
    BITFLIP_IND[95] <= 8'd95;
    BITFLIP_IND[96] <= 8'd96;
    BITFLIP_IND[97] <= 8'd97;
    BITFLIP_IND[98] <= 8'd98;
    BITFLIP_IND[99] <= 8'd99;
    BITFLIP_IND[100] <= 8'd100;
    BITFLIP_IND[101] <= 8'd101;
    BITFLIP_IND[102] <= 8'd102;
    BITFLIP_IND[103] <= 8'd103;
    BITFLIP_IND[104] <= 8'd104;
    BITFLIP_IND[105] <= 8'd105;
    BITFLIP_IND[106] <= 8'd106;
    BITFLIP_IND[107] <= 8'd107;
    BITFLIP_IND[108] <= 8'd108;
    BITFLIP_IND[109] <= 8'd109;
    BITFLIP_IND[110] <= 8'd110;
    BITFLIP_IND[111] <= 8'd111;
    BITFLIP_IND[112] <= 8'd112;
    BITFLIP_IND[113] <= 8'd113;
    BITFLIP_IND[114] <= 8'd114;
    BITFLIP_IND[115] <= 8'd115;
    BITFLIP_IND[116] <= 8'd116;
    BITFLIP_IND[117] <= 8'd117;
    BITFLIP_IND[118] <= 8'd118;
    BITFLIP_IND[119] <= 8'd119;
    BITFLIP_IND[120] <= 8'd120;
    BITFLIP_IND[121] <= 8'd121;
    BITFLIP_IND[122] <= 8'd122;
    BITFLIP_IND[123] <= 8'd123;
    BITFLIP_IND[124] <= 8'd124;
    BITFLIP_IND[125] <= 8'd125;
    BITFLIP_IND[126] <= 8'd126;
    BITFLIP_IND[127] <= 8'd127;
    BITFLIP_IND[128] <= 8'd128;
    BITFLIP_IND[129] <= 8'd129;
    BITFLIP_IND[130] <= 8'd130;
    BITFLIP_IND[131] <= 8'd131;
    BITFLIP_IND[132] <= 8'd132;
    BITFLIP_IND[133] <= 8'd133;
    BITFLIP_IND[134] <= 8'd134;
    BITFLIP_IND[135] <= 8'd135;
    BITFLIP_IND[136] <= 8'd136;
    BITFLIP_IND[137] <= 8'd137;
    BITFLIP_IND[138] <= 8'd138;
    BITFLIP_IND[139] <= 8'd139;
    BITFLIP_IND[140] <= 8'd140;
    BITFLIP_IND[141] <= 8'd141;
    BITFLIP_IND[142] <= 8'd142;
    BITFLIP_IND[143] <= 8'd143;
    BITFLIP_IND[144] <= 8'd144;
    BITFLIP_IND[145] <= 8'd145;
    BITFLIP_IND[146] <= 8'd146;
    BITFLIP_IND[147] <= 8'd147;
    BITFLIP_IND[148] <= 8'd148;
    BITFLIP_IND[149] <= 8'd149;
    BITFLIP_IND[150] <= 8'd150;
    BITFLIP_IND[151] <= 8'd151;
    BITFLIP_IND[152] <= 8'd152;
    BITFLIP_IND[153] <= 8'd153;
    BITFLIP_IND[154] <= 8'd154;
    BITFLIP_IND[155] <= 8'd155;
    BITFLIP_IND[156] <= 8'd156;
    BITFLIP_IND[157] <= 8'd157;
    BITFLIP_IND[158] <= 8'd158;
    BITFLIP_IND[159] <= 8'd159;
    BITFLIP_IND[160] <= 8'd160;
    BITFLIP_IND[161] <= 8'd161;
    BITFLIP_IND[162] <= 8'd162;
    BITFLIP_IND[163] <= 8'd163;
    BITFLIP_IND[164] <= 8'd164;
    BITFLIP_IND[165] <= 8'd165;
    BITFLIP_IND[166] <= 8'd166;
    BITFLIP_IND[167] <= 8'd167;
    BITFLIP_IND[168] <= 8'd168;
    BITFLIP_IND[169] <= 8'd169;
    BITFLIP_IND[170] <= 8'd170;
    BITFLIP_IND[171] <= 8'd171;
    BITFLIP_IND[172] <= 8'd172;
    BITFLIP_IND[173] <= 8'd173;
    BITFLIP_IND[174] <= 8'd174;
    BITFLIP_IND[175] <= 8'd175;
    BITFLIP_IND[176] <= 8'd176;
    BITFLIP_IND[177] <= 8'd177;
    BITFLIP_IND[178] <= 8'd178;
    BITFLIP_IND[179] <= 8'd179;
    BITFLIP_IND[180] <= 8'd180;
    BITFLIP_IND[181] <= 8'd181;
    BITFLIP_IND[182] <= 8'd182;
    BITFLIP_IND[183] <= 8'd183;
    BITFLIP_IND[184] <= 8'd184;
    BITFLIP_IND[185] <= 8'd185;
    BITFLIP_IND[186] <= 8'd186;
    BITFLIP_IND[187] <= 8'd187;
    BITFLIP_IND[188] <= 8'd188;
    BITFLIP_IND[189] <= 8'd189;
    BITFLIP_IND[190] <= 8'd190;
    BITFLIP_IND[191] <= 8'd191;
    BITFLIP_IND[192] <= 8'd192;
    BITFLIP_IND[193] <= 8'd193;
    BITFLIP_IND[194] <= 8'd194;
    BITFLIP_IND[195] <= 8'd195;
    BITFLIP_IND[196] <= 8'd196;
    BITFLIP_IND[197] <= 8'd197;
    BITFLIP_IND[198] <= 8'd198;
    BITFLIP_IND[199] <= 8'd199;
    BITFLIP_IND[200] <= 8'd200;
    BITFLIP_IND[201] <= 8'd201;
    BITFLIP_IND[202] <= 8'd202;
    BITFLIP_IND[203] <= 8'd203;
    BITFLIP_IND[204] <= 8'd204;
    BITFLIP_IND[205] <= 8'd205;
    BITFLIP_IND[206] <= 8'd206;
    BITFLIP_IND[207] <= 8'd207;
    BITFLIP_IND[208] <= 8'd208;
    BITFLIP_IND[209] <= 8'd209;
    BITFLIP_IND[210] <= 8'd210;
    BITFLIP_IND[211] <= 8'd211;
    BITFLIP_IND[212] <= 8'd212;
    BITFLIP_IND[213] <= 8'd213;
    BITFLIP_IND[214] <= 8'd214;
    BITFLIP_IND[215] <= 8'd215;
    BITFLIP_IND[216] <= 8'd216;
    BITFLIP_IND[217] <= 8'd217;
    BITFLIP_IND[218] <= 8'd218;
    BITFLIP_IND[219] <= 8'd219;
    BITFLIP_IND[220] <= 8'd220;
    BITFLIP_IND[221] <= 8'd221;
    BITFLIP_IND[222] <= 8'd222;
    BITFLIP_IND[223] <= 8'd223;
    BITFLIP_IND[224] <= 8'd224;
    BITFLIP_IND[225] <= 8'd225;
    BITFLIP_IND[226] <= 8'd226;
    BITFLIP_IND[227] <= 8'd227;
    BITFLIP_IND[228] <= 8'd228;
    BITFLIP_IND[229] <= 8'd229;
    BITFLIP_IND[230] <= 8'd230;
    BITFLIP_IND[231] <= 8'd231;
    BITFLIP_IND[232] <= 8'd232;
    BITFLIP_IND[233] <= 8'd233;
    BITFLIP_IND[234] <= 8'd234;
    BITFLIP_IND[235] <= 8'd235;
    BITFLIP_IND[236] <= 8'd236;
    BITFLIP_IND[237] <= 8'd237;
    BITFLIP_IND[238] <= 8'd238;
    BITFLIP_IND[239] <= 8'd239;
    BITFLIP_IND[240] <= 8'd240;
    BITFLIP_IND[241] <= 8'd241;
    BITFLIP_IND[242] <= 8'd242;
    BITFLIP_IND[243] <= 8'd243;
    BITFLIP_IND[244] <= 8'd244;
    BITFLIP_IND[245] <= 8'd245;
    BITFLIP_IND[246] <= 8'd246;
    BITFLIP_IND[247] <= 8'd247;
    BITFLIP_IND[248] <= 8'd248;
    BITFLIP_IND[249] <= 8'd249;
    BITFLIP_IND[250] <= 8'd250;
    BITFLIP_IND[251] <= 8'd251;
    BITFLIP_IND[252] <= 8'd252;
    BITFLIP_IND[253] <= 8'd253;
    BITFLIP_IND[254] <= 8'd254;
    BITFLIP_IND[255] <= 8'd255;
end

    // Stage FSM
    reg [3:0]state;
    //--------------------------- ila debug signals ------------------------
    assign state_fft = state;
    //----------------------------------------------------------------------
    localparam IDLE = 4'b0000, STAGE1 = 4'b0001, STAGE2 = 4'b0010, STAGE3 = 4'b0011, STAGE4 = 4'b0100, STAGE5 = 4'b0101, STAGE6 = 4'b0110, STAGE7 = 4'b0111, STAGE8 = 4'b1000, BIT_FLIP_STAGE = 4'b1001, CLEANUP = 4'b1010;
    reg [8:0]st_ctr;
    reg [2:0]flipper;
    reg latency_ctrl; // to tackle the 1 cycle latency caused on ram address setting
    reg [((2*WIDTH)-1):0] d1, d2;
    reg [WIDTH-1 : 0] d1_1, d1_2, d2_1, d2_2;
    always@(posedge clk or negedge rst) begin
        if(rst == 1'b0) begin
            w_real <= 0;
            w_imag <= 0;
            in1_real <= 0;
            in1_imag <= 0;
            in2_real <=0;
            in2_imag <= 0;
            st_ctr <= 4'b0;
            flipper <= 1'b0;
            addr_tw <= 0;
            done <= 1'b0;
            addrb <= 0;
            addra <= 0;
            douta <= 0;
            state <= IDLE;
            wr <= 0;
            tw<=0;
            latency_ctrl <= 0;
            d_fifo_ram <= 0;
            wr_fifo_ram <= 0;
            addr_fifo_ram <= 0;
            d1 <= 0;
            d2 <= 0;
            d2_1 <= 0;
            d2_2 <= 0;
            d1_1 <= 0;
            d1_2 <= 0;
        end else begin
            case(state)
                IDLE : begin
                    done <= 1'b0;
                    wr <= 0;
                    if(trig) begin 
                        state <= STAGE1;
                    end 
                end
                STAGE1 : begin
                    if(st_ctr > 255) begin
                        state <= STAGE2;
                        addrb <= 0;
                        addra <= 0;
                        st_ctr <= 0;
                        flipper <= 0;
                        wr <= 0;
                        latency_ctrl <= 0;
                    end else begin
                        if(flipper == 0 || flipper == 2) begin
                            // sample fetch
                            wr <= 0;
                            addrb <= STAGE1_IND[st_ctr];
                            if(latency_ctrl) begin
                                flipper <= flipper + 1;
                            end
                            if(flipper == 2 && latency_ctrl) begin
                                // twiddle factor fetch
                                tw <= dout_tw;
                                addr_tw <= addr_tw + 1;
                            end
                            latency_ctrl <= latency_ctrl + 1;
                        end else if(flipper == 1) begin
                                in1_real<= doutb[(WIDTH - 1) : 0];     
                                in1_imag<= doutb[((2*WIDTH) - 1) : WIDTH];
                                flipper <= flipper + 1;
                                st_ctr <= st_ctr + 1;
                            end else if(flipper == 3) begin
                                in2_real<= doutb[WIDTH - 1 : 0];
                                in2_imag<= doutb[2*WIDTH - 1 : WIDTH];
                                flipper <= flipper + 1;
                                w_real <= {{8{tw[11]}}, tw[11:0]};
                                w_imag <= {{8{tw[23]}}, tw[23:12]};
                        end else if(flipper == 4) begin
                            douta <= {out1_imag, out1_real};
                            wr <= 1'b1;
                            flipper <= flipper + 1;
                            addra <= STAGE1_IND[st_ctr - 1];
                        end else if(flipper == 5) begin
                            wr <= 1'b1;
                            douta <= {out2_imag, out2_real};
                            flipper <= 0;
                            addra <= STAGE1_IND[st_ctr];
                            st_ctr <= st_ctr + 1;
                        end
                    end
                end
                STAGE2 : begin
                    if(st_ctr > 255) begin
                        state <= STAGE3;
                        addrb <= 0;
                        addra <= 0;
                        st_ctr <= 0;
                        flipper <= 0;
                        wr <= 0;
                        latency_ctrl <= 0;
                    end else begin
                        if(flipper == 0 || flipper == 2) begin
                            wr <= 0;
                            // sample fetch
                            addrb <= STAGE2_IND[st_ctr];
                            if(latency_ctrl) begin
                                flipper <= flipper + 1;
                            end
                            if(flipper == 2 && latency_ctrl) begin
                                // twiddle factor fetch
                                tw <= dout_tw;
                                addr_tw <= addr_tw + 1;
                            end
                            latency_ctrl <= latency_ctrl + 1;
                        end else if(flipper == 1) begin
                                in1_real<= doutb[WIDTH - 1 : 0];       
                                in1_imag<= doutb[2*WIDTH - 1 : WIDTH]; 
                                flipper <= flipper + 1;
                                st_ctr <= st_ctr + 1;
                            end else if(flipper == 3) begin
                                in2_real<= doutb[WIDTH - 1 : 0];       
                                in2_imag<= doutb[2*WIDTH - 1 : WIDTH]; 
                                w_real <= {{8{tw[11]}}, tw[11:0]}; 
                                w_imag <= {{8{tw[23]}}, tw[23:12]};
                                flipper <= flipper + 1;
                        end else if(flipper == 4) begin
                            douta <= {out1_imag, out1_real};
                            flipper <= flipper + 1;
                            addra <= STAGE2_IND[st_ctr - 1];
                            wr <= 1'b1;
                        end else if(flipper == 5) begin
                            douta <= {out2_imag, out2_real};
                            flipper <= 0;
                            addra <= STAGE2_IND[st_ctr]; 
                            st_ctr <= st_ctr + 1;
                            wr <= 1'b1;
                        end
                    end
                end
                
                STAGE3 : begin
                    if(st_ctr > 255) begin
                        state <= STAGE4;
                        addrb <= 0;
                        addra <= 0;
                        st_ctr <= 0;
                        flipper <= 0;
                        wr <= 0;
                        latency_ctrl <= 0;
                    end else begin
                        if(flipper == 0 || flipper == 2) begin
                            wr <= 0;
                            // sample fetch
                            addrb <= STAGE3_IND[st_ctr];
                            if(latency_ctrl) begin
                                flipper <= flipper + 1;
                            end
                            if(flipper == 2 && latency_ctrl) begin
                                // twiddle factor fetch
                                tw <= dout_tw;
                                addr_tw <= addr_tw + 1;
                            end
                            latency_ctrl <= latency_ctrl + 1;
                        end else if(flipper == 1) begin
                                in1_real<= doutb[WIDTH - 1 : 0];       
                                in1_imag<= doutb[2*WIDTH - 1 : WIDTH]; 
                                flipper <= flipper + 1;
                                st_ctr <= st_ctr + 1;
                            end else if(flipper == 3) begin
                                in2_real<= doutb[WIDTH - 1 : 0];       
                                in2_imag<= doutb[2*WIDTH - 1 : WIDTH]; 
                                w_real <= {{8{tw[11]}}, tw[11:0]}; 
                                w_imag <= {{8{tw[23]}}, tw[23:12]};
                                flipper <= flipper + 1;
                        end else if(flipper == 4) begin
                            douta <= {out1_imag, out1_real};
                            flipper <= flipper + 1;
                            addra <= STAGE3_IND[st_ctr - 1];
                            wr <= 1'b1;
                        end else if(flipper == 5) begin
                            douta <= {out2_imag, out2_real};
                            flipper <= 0;
                            addra <= STAGE3_IND[st_ctr]; 
                            st_ctr <= st_ctr + 1;
                            wr <= 1'b1;
                        end
                    end
                end
                
                STAGE4 : begin
                    if(st_ctr > 255) begin
                        state <= STAGE5;
                        addrb <= 0;
                        addra <= 0;
                        st_ctr <= 0;
                        flipper <= 0;
                        wr <= 0;
                        latency_ctrl <= 0;
                    end else begin
                        if(flipper == 0 || flipper == 2) begin
                            wr <= 0;
                            // sample fetch
                            addrb <= STAGE4_IND[st_ctr];
                            if(latency_ctrl) begin
                                flipper <= flipper + 1;
                            end
                            if(flipper == 2 && latency_ctrl) begin
                                // twiddle factor fetch
                                tw <= dout_tw;
                                addr_tw <= addr_tw + 1;
                            end
                            latency_ctrl <= latency_ctrl + 1;
                        end else if(flipper == 1) begin
                                in1_real<= doutb[WIDTH - 1 : 0];       
                                in1_imag<= doutb[2*WIDTH - 1 : WIDTH]; 
                                flipper <= flipper + 1;
                                st_ctr <= st_ctr + 1;
                            end else if(flipper == 3) begin
                                in2_real<= doutb[WIDTH - 1 : 0];       
                                in2_imag<= doutb[2*WIDTH - 1 : WIDTH]; 
                                w_real <= {{8{tw[11]}}, tw[11:0]}; 
                                w_imag <= {{8{tw[23]}}, tw[23:12]};
                                flipper <= flipper + 1;
                        end else if(flipper == 4) begin
                            douta <= {out1_imag, out1_real};
                            flipper <= flipper + 1;
                            addra <= STAGE4_IND[st_ctr - 1];
                            wr <= 1'b1;
                        end else if(flipper == 5) begin
                            douta <= {out2_imag, out2_real};
                            flipper <= 0;
                            addra <= STAGE4_IND[st_ctr]; 
                            st_ctr <= st_ctr + 1;
                            wr <= 1'b1;
                        end
                    end
                end
                
                STAGE5 : begin
                    if(st_ctr > 255) begin
                        state <= STAGE6;
                        addrb <= 0;
                        addra <= 0;
                        st_ctr <= 0;
                        flipper <= 0;
                        wr <= 0;
                        latency_ctrl <= 0;
                    end else begin
                        if(flipper == 0 || flipper == 2) begin
                            wr <= 0;
                            // sample fetch
                            addrb <= STAGE5_IND[st_ctr];
                            if(latency_ctrl) begin
                                flipper <= flipper + 1;
                            end
                            if(flipper == 2 && latency_ctrl) begin
                                // twiddle factor fetch
                                tw <= dout_tw;
                                addr_tw <= addr_tw + 1;
                            end
                            latency_ctrl <= latency_ctrl + 1;
                        end else if(flipper == 1) begin
                                in1_real<= doutb[WIDTH - 1 : 0];       
                                in1_imag<= doutb[2*WIDTH - 1 : WIDTH]; 
                                flipper <= flipper + 1;
                                st_ctr <= st_ctr + 1;
                            end else if(flipper == 3) begin
                                in2_real<= doutb[WIDTH - 1 : 0];       
                                in2_imag<= doutb[2*WIDTH - 1 : WIDTH]; 
                                w_real <= {{8{tw[11]}}, tw[11:0]}; 
                                w_imag <= {{8{tw[23]}}, tw[23:12]};
                                flipper <= flipper + 1;
                        end else if(flipper == 4) begin
                            douta <= {out1_imag, out1_real};
                            flipper <= flipper + 1;
                            addra <= STAGE5_IND[st_ctr - 1];
                            wr <= 1'b1;
                        end else if(flipper == 5) begin
                            douta <= {out2_imag, out2_real};
                            flipper <= 0;
                            addra <= STAGE5_IND[st_ctr]; 
                            st_ctr <= st_ctr + 1;
                            wr <= 1'b1;
                        end
                    end
                end
                
                STAGE6 : begin
                    if(st_ctr > 255) begin
                        state <= STAGE7;
                        addrb <= 0;
                        addra <= 0;
                        st_ctr <= 0;
                        flipper <= 0;
                        wr <= 0;
                        latency_ctrl <= 0;
                    end else begin
                        if(flipper == 0 || flipper == 2) begin
                            wr <= 0;
                            // sample fetch
                            addrb <= STAGE6_IND[st_ctr];
                            if(latency_ctrl) begin
                                flipper <= flipper + 1;
                            end
                            if(flipper == 2 && latency_ctrl) begin
                                // twiddle factor fetch
                                tw <= dout_tw;
                                addr_tw <= addr_tw + 1;
                            end
                            latency_ctrl <= latency_ctrl + 1;
                        end else if(flipper == 1) begin
                                in1_real<= doutb[WIDTH - 1 : 0];       
                                in1_imag<= doutb[2*WIDTH - 1 : WIDTH]; 
                                flipper <= flipper + 1;
                                st_ctr <= st_ctr + 1;
                            end else if(flipper == 3) begin
                                in2_real<= doutb[WIDTH - 1 : 0];       
                                in2_imag<= doutb[2*WIDTH - 1 : WIDTH]; 
                                w_real <= {{8{tw[11]}}, tw[11:0]}; 
                                w_imag <= {{8{tw[23]}}, tw[23:12]};
                                flipper <= flipper + 1;
                        end else if(flipper == 4) begin
                            douta <= {out1_imag, out1_real};
                            flipper <= flipper + 1;
                            addra <= STAGE6_IND[st_ctr - 1];
                            wr <= 1'b1;
                        end else if(flipper == 5) begin
                            douta <= {out2_imag, out2_real};
                            flipper <= 0;
                            addra <= STAGE6_IND[st_ctr]; 
                            st_ctr <= st_ctr + 1;
                            wr <= 1'b1;
                        end
                    end
                end
                
                STAGE7 : begin
                    if(st_ctr > 255) begin
                        state <= STAGE8;
                        addrb <= 0;
                        addra <= 0;
                        st_ctr <= 0;
                        flipper <= 0;
                        wr <= 0;
                        latency_ctrl <= 0;
                    end else begin
                        if(flipper == 0 || flipper == 2) begin
                            wr <= 0;
                            // sample fetch
                            addrb <= STAGE7_IND[st_ctr];
                            if(latency_ctrl) begin
                                flipper <= flipper + 1;
                            end
                            if(flipper == 2 && latency_ctrl) begin
                                // twiddle factor fetch
                                tw <= dout_tw;
                                addr_tw <= addr_tw + 1;
                            end
                            latency_ctrl <= latency_ctrl + 1;
                        end else if(flipper == 1) begin
                                in1_real<= doutb[WIDTH - 1 : 0];       
                                in1_imag<= doutb[2*WIDTH - 1 : WIDTH]; 
                                flipper <= flipper + 1;
                                st_ctr <= st_ctr + 1;
                            end else if(flipper == 3) begin
                                in2_real<= doutb[WIDTH - 1 : 0];       
                                in2_imag<= doutb[2*WIDTH - 1 : WIDTH]; 
                                w_real <= {{8{tw[11]}}, tw[11:0]}; 
                                w_imag <= {{8{tw[23]}}, tw[23:12]};
                                flipper <= flipper + 1;
                        end else if(flipper == 4) begin
                            douta <= {out1_imag, out1_real};
                            flipper <= flipper + 1;
                            addra <= STAGE7_IND[st_ctr - 1];
                            wr <= 1'b1;
                        end else if(flipper == 5) begin
                            douta <= {out2_imag, out2_real};
                            flipper <= 0;
                            addra <= STAGE7_IND[st_ctr]; 
                            st_ctr <= st_ctr + 1;
                            wr <= 1'b1;
                        end
                    end
                end
                
                STAGE8 : begin  // LAST STAGE OF FFT 
                    if(st_ctr > 255) begin
                        state <= BIT_FLIP_STAGE;
                        addrb <= 0;
                        addra <= 0;
                        st_ctr <= 0;
                        addr_tw <= 0;
                        flipper <= 0;
                        done <= 1'b0;
                        wr <= 0;
                        latency_ctrl <= 0;
                    end else begin
                        if(flipper == 0 || flipper == 2) begin
                            wr <= 0;
                            // sample fetch
                            addrb <= STAGE8_IND[st_ctr];
                            if(latency_ctrl) begin
                                flipper <= flipper + 1;
                            end
                            if(flipper == 2 && latency_ctrl) begin
                                // twiddle factor fetch
                                tw <= dout_tw;
                                addr_tw <= addr_tw + 1;
                            end
                            latency_ctrl <= latency_ctrl + 1;
                        end else if(flipper == 1) begin
                                in1_real<= doutb[WIDTH - 1 : 0];       
                                in1_imag<= doutb[2*WIDTH - 1 : WIDTH]; 
                                flipper <= flipper + 1;
                                st_ctr <= st_ctr + 1;
                            end else if(flipper == 3) begin
                                in2_real<= doutb[WIDTH - 1 : 0];       
                                in2_imag<= doutb[2*WIDTH - 1 : WIDTH]; 
                                w_real <= {{8{tw[11]}}, tw[11:0]}; 
                                w_imag <= {{8{tw[23]}}, tw[23:12]};
                                flipper <= flipper + 1;
                        end else if(flipper == 4) begin
                            douta <= {out1_imag, out1_real};
                            flipper <= flipper + 1;
                            addra <= STAGE8_IND[st_ctr - 1];
                            wr <= 1'b1;
                        end else if(flipper == 5) begin
                            douta <= {out2_imag, out2_real};
                            flipper <= 0;
                            addra <= STAGE8_IND[st_ctr];
                            st_ctr <= st_ctr + 1;
                            wr <= 1'b1;
                        end
                    end
                end
                BIT_FLIP_STAGE : begin
                    if(st_ctr > 255) begin
                        state <= CLEANUP;
                        addrb <= 0;
                        addra <= 0;
                        st_ctr <= 0;
                        flipper <= 0;
                        wr_fifo_ram <= 0;
                        latency_ctrl <= 0;
                        done <= 1'b1;
                    end else begin
                        if(flipper == 0 || flipper == 2) begin
                            // sample fetch
                            wr_fifo_ram <= 0;
                            addrb <= BITFLIP_IND[st_ctr]; 
                            
                            if(latency_ctrl) begin
                                flipper <= flipper + 1;
                            end          
                            
                            latency_ctrl <= latency_ctrl + 1;
                        end else if(flipper == 1) begin
                                d1 <= doutb;
                                flipper <= flipper + 1;
                                st_ctr <= st_ctr + 1;
                            end else if(flipper == 3) begin
                                d2 <= doutb;
                                flipper <= flipper + 1;
                        end else if(flipper == 4) begin
                            d1_1 = ((d1[2*WIDTH - 1 : WIDTH])>>>SHIFT_FACTOR);
                            d1_2 = ((d1[WIDTH - 1 : 0])>>>SHIFT_FACTOR);
                            d_fifo_ram <= {d1_1[11:0], d1_2[11:0]};
//                            d_fifo_ram <= 24'hffffff;  // for debug
                            wr_fifo_ram <= 1'b1;
                            flipper <= flipper + 1;
                            addr_fifo_ram <= {STAGE1_IND[st_ctr - 1], 2'b0};
                        end else if(flipper == 5) begin
                            wr_fifo_ram <= 1'b1;
                            d2_1 = ((d2[2*WIDTH - 1 : WIDTH])>>>SHIFT_FACTOR);
                            d2_2 = ((d2[WIDTH - 1 : 0])>>>SHIFT_FACTOR);  
                            d_fifo_ram <=  {d2_1[11:0], d2_2[11:0]};
//                            d_fifo_ram <= 24'hffffff;  // for debug
                            flipper <= 0;
                            addr_fifo_ram <= {STAGE1_IND[st_ctr], 2'b0};
                            st_ctr <= st_ctr + 1;
                        end
                    end
                end
                
                CLEANUP : begin
                    w_real <= 0;
                    w_imag <= 0;
                    in1_real <= 0;
                    in1_imag <= 0;
                    in2_real <=0;
                    in2_imag <= 0;
                    st_ctr <= 4'b0;
                    flipper <= 1'b0;
                    addr_tw <= 1'b0;
                    done <= 1'b1;
                    addrb <= 0;
                    addra <= 0;
                    douta <= 0;
                    state <= IDLE;
                    wr <= 0;
                    tw<=0;
                    latency_ctrl <= 0;
                    d_fifo_ram <= 0;
                    wr_fifo_ram <= 0;
                    addr_fifo_ram <= 0;
                    d1 <= 0;
                    d2 <= 0;
                end
            endcase
        end
    end
    
    
endmodule
